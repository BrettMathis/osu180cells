module ffra (clk,
    rst,
    vdd,
    vss,
    a,
    b,
    ci,
    o);
 input clk;
 input rst;
 input vdd;
 input vss;
 input [7:0] a;
 input [7:0] b;
 input [15:0] ci;
 output [15:0] o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire \o_tmp[0][0] ;
 wire \o_tmp[0][10] ;
 wire \o_tmp[0][11] ;
 wire \o_tmp[0][12] ;
 wire \o_tmp[0][13] ;
 wire \o_tmp[0][14] ;
 wire \o_tmp[0][15] ;
 wire \o_tmp[0][1] ;
 wire \o_tmp[0][2] ;
 wire \o_tmp[0][3] ;
 wire \o_tmp[0][4] ;
 wire \o_tmp[0][5] ;
 wire \o_tmp[0][6] ;
 wire \o_tmp[0][7] ;
 wire \o_tmp[0][8] ;
 wire \o_tmp[0][9] ;
 wire \o_tmp[1][0] ;
 wire \o_tmp[1][10] ;
 wire \o_tmp[1][11] ;
 wire \o_tmp[1][12] ;
 wire \o_tmp[1][13] ;
 wire \o_tmp[1][14] ;
 wire \o_tmp[1][15] ;
 wire \o_tmp[1][1] ;
 wire \o_tmp[1][2] ;
 wire \o_tmp[1][3] ;
 wire \o_tmp[1][4] ;
 wire \o_tmp[1][5] ;
 wire \o_tmp[1][6] ;
 wire \o_tmp[1][7] ;
 wire \o_tmp[1][8] ;
 wire \o_tmp[1][9] ;
 wire \o_tmp[2][0] ;
 wire \o_tmp[2][10] ;
 wire \o_tmp[2][11] ;
 wire \o_tmp[2][12] ;
 wire \o_tmp[2][13] ;
 wire \o_tmp[2][14] ;
 wire \o_tmp[2][15] ;
 wire \o_tmp[2][1] ;
 wire \o_tmp[2][2] ;
 wire \o_tmp[2][3] ;
 wire \o_tmp[2][4] ;
 wire \o_tmp[2][5] ;
 wire \o_tmp[2][6] ;
 wire \o_tmp[2][7] ;
 wire \o_tmp[2][8] ;
 wire \o_tmp[2][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;

 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0522_ (.VDD(vdd),
    .VSS(vss),
    .A(net9),
    .Y(_0405_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0523_ (.VDD(vdd),
    .VSS(vss),
    .A(_0405_),
    .Y(_0411_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0524_ (.VDD(vdd),
    .VSS(vss),
    .A(net1),
    .Y(_0412_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0525_ (.VDD(vdd),
    .VSS(vss),
    .A(_0412_),
    .Y(_0413_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0526_ (.VDD(vdd),
    .VSS(vss),
    .A(_0411_),
    .B(_0413_),
    .Y(_0414_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0527_ (.VDD(vdd),
    .VSS(vss),
    .A(net17),
    .B(_0414_),
    .Y(_0415_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0528_ (.VDD(vdd),
    .VSS(vss),
    .A(_0415_),
    .Y(_0000_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0529_ (.VDD(vdd),
    .VSS(vss),
    .A(net17),
    .Y(_0416_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0530_ (.VDD(vdd),
    .VSS(vss),
    .A(_0416_),
    .B(_0414_),
    .Y(_0417_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0531_ (.VDD(vdd),
    .VSS(vss),
    .A(net10),
    .Y(_0418_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0532_ (.VDD(vdd),
    .VSS(vss),
    .A(_0418_),
    .Y(_0419_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0533_ (.VDD(vdd),
    .VSS(vss),
    .A(_0419_),
    .B(_0413_),
    .Y(_0420_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0534_ (.VDD(vdd),
    .VSS(vss),
    .A(net2),
    .Y(_0421_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0535_ (.VDD(vdd),
    .VSS(vss),
    .A(_0421_),
    .Y(_0422_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0536_ (.VDD(vdd),
    .VSS(vss),
    .A(_0422_),
    .B(_0411_),
    .Y(_0423_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0537_ (.VDD(vdd),
    .VSS(vss),
    .A(net24),
    .B(_0423_),
    .Y(_0424_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0538_ (.VDD(vdd),
    .VSS(vss),
    .A(_0420_),
    .B(_0424_),
    .Y(_0425_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0539_ (.VDD(vdd),
    .VSS(vss),
    .A(_0417_),
    .B(_0425_),
    .Y(_0426_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0540_ (.VDD(vdd),
    .VSS(vss),
    .A(_0426_),
    .Y(_0427_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0541_ (.VDD(vdd),
    .VSS(vss),
    .A(_0417_),
    .B(_0425_),
    .Y(_0428_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0542_ (.VDD(vdd),
    .VSS(vss),
    .A(_0427_),
    .B(_0428_),
    .Y(_0429_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0543_ (.VDD(vdd),
    .VSS(vss),
    .A(_0429_),
    .Y(_0001_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0544_ (.VDD(vdd),
    .VSS(vss),
    .A(net11),
    .Y(_0430_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0545_ (.VDD(vdd),
    .VSS(vss),
    .A(net1),
    .B(_0430_),
    .Y(_0431_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0546_ (.VDD(vdd),
    .VSS(vss),
    .A(_0421_),
    .B(_0419_),
    .Y(_0432_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0547_ (.VDD(vdd),
    .VSS(vss),
    .A(net3),
    .Y(_0433_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0548_ (.VDD(vdd),
    .VSS(vss),
    .A(_0411_),
    .B(_0433_),
    .Y(_0434_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0549_ (.VDD(vdd),
    .VSS(vss),
    .A(net25),
    .B(_0434_),
    .Y(_0435_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0550_ (.VDD(vdd),
    .VSS(vss),
    .A(_0432_),
    .B(_0435_),
    .Y(_0436_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0551_ (.VDD(vdd),
    .VSS(vss),
    .A(net24),
    .B(_0423_),
    .Y(_0437_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0552_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0420_),
    .A1(_0424_),
    .B(_0437_),
    .Y(_0438_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0553_ (.VDD(vdd),
    .VSS(vss),
    .A(_0436_),
    .B(_0438_),
    .Y(_0439_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0554_ (.VDD(vdd),
    .VSS(vss),
    .A(_0431_),
    .B(_0439_),
    .Y(_0440_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0555_ (.VDD(vdd),
    .VSS(vss),
    .A(_0426_),
    .B(_0440_),
    .Y(_0441_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0556_ (.VDD(vdd),
    .VSS(vss),
    .A(_0441_),
    .Y(_0002_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0557_ (.VDD(vdd),
    .VSS(vss),
    .A(_0427_),
    .B(_0440_),
    .Y(_0442_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0558_ (.VDD(vdd),
    .VSS(vss),
    .A(_0436_),
    .B(_0438_),
    .Y(_0443_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0559_ (.VDD(vdd),
    .VSS(vss),
    .A(_0436_),
    .B(_0438_),
    .Y(_0444_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0560_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0431_),
    .A1(_0443_),
    .B(_0444_),
    .Y(_0445_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0561_ (.VDD(vdd),
    .VSS(vss),
    .A(net12),
    .Y(_0446_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0562_ (.VDD(vdd),
    .VSS(vss),
    .A(_0421_),
    .B(_0446_),
    .Y(_0447_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0563_ (.VDD(vdd),
    .VSS(vss),
    .A(_0431_),
    .B(_0447_),
    .Y(_0448_));
 gf180mcu_osu_sc_gp9t3v3__aoi22_1 _0564_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0422_),
    .A1(_0430_),
    .B0(_0446_),
    .B1(_0412_),
    .Y(_0449_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0565_ (.VDD(vdd),
    .VSS(vss),
    .A(_0448_),
    .B(_0449_),
    .Y(_0450_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0566_ (.VDD(vdd),
    .VSS(vss),
    .A(net3),
    .Y(_0451_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0567_ (.VDD(vdd),
    .VSS(vss),
    .A(_0419_),
    .B(_0451_),
    .Y(_0452_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0568_ (.VDD(vdd),
    .VSS(vss),
    .A(net4),
    .Y(_0453_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0569_ (.VDD(vdd),
    .VSS(vss),
    .A(_0411_),
    .B(_0453_),
    .Y(_0454_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0570_ (.VDD(vdd),
    .VSS(vss),
    .A(net26),
    .B(_0454_),
    .Y(_0455_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0571_ (.VDD(vdd),
    .VSS(vss),
    .A(_0452_),
    .B(_0455_),
    .Y(_0456_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0572_ (.VDD(vdd),
    .VSS(vss),
    .A(net25),
    .B(_0434_),
    .Y(_0457_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0573_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0432_),
    .A1(_0435_),
    .B(_0457_),
    .Y(_0016_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0574_ (.VDD(vdd),
    .VSS(vss),
    .A(_0456_),
    .B(_0016_),
    .Y(_0017_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0575_ (.VDD(vdd),
    .VSS(vss),
    .A(_0450_),
    .B(_0017_),
    .Y(_0018_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0576_ (.VDD(vdd),
    .VSS(vss),
    .A(_0445_),
    .B(_0018_),
    .Y(_0019_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0577_ (.VDD(vdd),
    .VSS(vss),
    .A(_0442_),
    .B(_0019_),
    .Y(_0020_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0578_ (.VDD(vdd),
    .VSS(vss),
    .A(_0020_),
    .Y(_0003_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0579_ (.VDD(vdd),
    .VSS(vss),
    .A(_0445_),
    .B(_0018_),
    .Y(_0021_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0580_ (.VDD(vdd),
    .VSS(vss),
    .A(_0021_),
    .Y(_0022_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0581_ (.VDD(vdd),
    .VSS(vss),
    .A(_0450_),
    .Y(_0023_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0582_ (.VDD(vdd),
    .VSS(vss),
    .A(_0456_),
    .B(_0016_),
    .Y(_0024_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0583_ (.VDD(vdd),
    .VSS(vss),
    .A(_0456_),
    .B(_0016_),
    .Y(_0025_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0584_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0023_),
    .A1(_0024_),
    .B(_0025_),
    .Y(_0026_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0585_ (.VDD(vdd),
    .VSS(vss),
    .A(net26),
    .B(_0454_),
    .Y(_0027_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0586_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0452_),
    .A1(_0455_),
    .B(_0027_),
    .Y(_0028_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0587_ (.VDD(vdd),
    .VSS(vss),
    .A(_0418_),
    .B(_0453_),
    .Y(_0029_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0588_ (.VDD(vdd),
    .VSS(vss),
    .A(_0405_),
    .B(net5),
    .Y(_0030_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0589_ (.VDD(vdd),
    .VSS(vss),
    .A(net27),
    .B(_0030_),
    .Y(_0031_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0590_ (.VDD(vdd),
    .VSS(vss),
    .A(_0029_),
    .B(_0031_),
    .Y(_0032_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0591_ (.VDD(vdd),
    .VSS(vss),
    .A(_0028_),
    .B(_0032_),
    .Y(_0033_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0592_ (.VDD(vdd),
    .VSS(vss),
    .A(net13),
    .Y(_0034_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0593_ (.VDD(vdd),
    .VSS(vss),
    .A(_0412_),
    .B(_0034_),
    .Y(_0035_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0594_ (.VDD(vdd),
    .VSS(vss),
    .A(_0433_),
    .B(_0430_),
    .Y(_0036_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0595_ (.VDD(vdd),
    .VSS(vss),
    .A(_0447_),
    .B(_0036_),
    .Y(_0037_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0596_ (.VDD(vdd),
    .VSS(vss),
    .A(_0035_),
    .B(_0037_),
    .Y(_0038_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0597_ (.VDD(vdd),
    .VSS(vss),
    .A(_0033_),
    .B(_0038_),
    .Y(_0039_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0598_ (.VDD(vdd),
    .VSS(vss),
    .A(_0026_),
    .B(_0039_),
    .Y(_0040_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0599_ (.VDD(vdd),
    .VSS(vss),
    .A(_0448_),
    .B(_0040_),
    .Y(_0041_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0600_ (.VDD(vdd),
    .VSS(vss),
    .A(_0022_),
    .B(_0041_),
    .Y(_0042_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0601_ (.VDD(vdd),
    .VSS(vss),
    .A(_0447_),
    .B(_0036_),
    .Y(_0043_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0602_ (.VDD(vdd),
    .VSS(vss),
    .A(_0035_),
    .B(_0037_),
    .Y(_0044_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0603_ (.VDD(vdd),
    .VSS(vss),
    .A(_0043_),
    .B(_0044_),
    .Y(_0045_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0604_ (.VDD(vdd),
    .VSS(vss),
    .A(net14),
    .Y(_0046_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0605_ (.VDD(vdd),
    .VSS(vss),
    .A(_0046_),
    .Y(_0047_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0606_ (.VDD(vdd),
    .VSS(vss),
    .A(_0413_),
    .B(_0047_),
    .Y(_0048_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0607_ (.VDD(vdd),
    .VSS(vss),
    .A(_0045_),
    .B(_0048_),
    .Y(_0049_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0608_ (.VDD(vdd),
    .VSS(vss),
    .A(_0045_),
    .B(_0048_),
    .Y(_0050_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0609_ (.VDD(vdd),
    .VSS(vss),
    .A(_0049_),
    .B(_0050_),
    .Y(_0051_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0610_ (.VDD(vdd),
    .VSS(vss),
    .A(net5),
    .Y(_0052_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0611_ (.VDD(vdd),
    .VSS(vss),
    .A(_0418_),
    .B(_0052_),
    .Y(_0053_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0612_ (.VDD(vdd),
    .VSS(vss),
    .A(_0405_),
    .B(net6),
    .Y(_0054_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0613_ (.VDD(vdd),
    .VSS(vss),
    .A(net28),
    .B(_0054_),
    .Y(_0055_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0614_ (.VDD(vdd),
    .VSS(vss),
    .A(_0053_),
    .B(_0055_),
    .Y(_0056_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0615_ (.VDD(vdd),
    .VSS(vss),
    .A(net27),
    .B(_0030_),
    .Y(_0057_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0616_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0029_),
    .A1(_0031_),
    .B(_0057_),
    .Y(_0058_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0617_ (.VDD(vdd),
    .VSS(vss),
    .A(_0056_),
    .B(_0058_),
    .Y(_0059_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0618_ (.VDD(vdd),
    .VSS(vss),
    .A(net13),
    .Y(_0060_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0619_ (.VDD(vdd),
    .VSS(vss),
    .A(_0421_),
    .B(_0060_),
    .Y(_0061_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0620_ (.VDD(vdd),
    .VSS(vss),
    .A(_0433_),
    .B(_0446_),
    .Y(_0062_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0621_ (.VDD(vdd),
    .VSS(vss),
    .A(net11),
    .Y(_0063_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0622_ (.VDD(vdd),
    .VSS(vss),
    .A(_0063_),
    .B(_0453_),
    .Y(_0064_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0623_ (.VDD(vdd),
    .VSS(vss),
    .A(_0062_),
    .B(_0064_),
    .Y(_0065_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0624_ (.VDD(vdd),
    .VSS(vss),
    .A(_0061_),
    .B(_0065_),
    .Y(_0066_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0625_ (.VDD(vdd),
    .VSS(vss),
    .A(_0059_),
    .B(_0066_),
    .Y(_0067_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0626_ (.VDD(vdd),
    .VSS(vss),
    .A(_0028_),
    .B(_0032_),
    .Y(_0068_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0627_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0033_),
    .A1(_0038_),
    .B(_0068_),
    .Y(_0069_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0628_ (.VDD(vdd),
    .VSS(vss),
    .A(_0067_),
    .B(_0069_),
    .Y(_0070_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0629_ (.VDD(vdd),
    .VSS(vss),
    .A(_0051_),
    .B(_0070_),
    .Y(_0071_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0630_ (.VDD(vdd),
    .VSS(vss),
    .A(_0026_),
    .B(_0039_),
    .Y(_0072_));
 gf180mcu_osu_sc_gp9t3v3__oai31_1 _0631_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0431_),
    .A1(_0447_),
    .A2(_0040_),
    .B(_0072_),
    .Y(_0073_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0632_ (.VDD(vdd),
    .VSS(vss),
    .A(_0071_),
    .B(_0073_),
    .Y(_0074_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0633_ (.VDD(vdd),
    .VSS(vss),
    .A(_0042_),
    .B(_0074_),
    .Y(_0075_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0634_ (.VDD(vdd),
    .VSS(vss),
    .A(_0442_),
    .B(_0019_),
    .Y(_0076_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0635_ (.VDD(vdd),
    .VSS(vss),
    .A(_0076_),
    .B(_0041_),
    .Y(_0077_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0636_ (.VDD(vdd),
    .VSS(vss),
    .A(_0075_),
    .B(_0077_),
    .Y(_0078_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0637_ (.VDD(vdd),
    .VSS(vss),
    .A(_0078_),
    .Y(_0011_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0638_ (.VDD(vdd),
    .VSS(vss),
    .A(_0071_),
    .Y(_0079_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0639_ (.VDD(vdd),
    .VSS(vss),
    .A(_0079_),
    .B(_0073_),
    .Y(_0080_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0640_ (.VDD(vdd),
    .VSS(vss),
    .A(net12),
    .Y(_0081_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0641_ (.VDD(vdd),
    .VSS(vss),
    .A(_0453_),
    .B(_0081_),
    .Y(_0082_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0642_ (.VDD(vdd),
    .VSS(vss),
    .A(_0036_),
    .B(_0082_),
    .Y(_0083_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0643_ (.VDD(vdd),
    .VSS(vss),
    .A(_0061_),
    .B(_0065_),
    .Y(_0084_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0644_ (.VDD(vdd),
    .VSS(vss),
    .A(_0083_),
    .B(_0084_),
    .Y(_0085_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0645_ (.VDD(vdd),
    .VSS(vss),
    .A(net2),
    .B(net15),
    .Y(_0086_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0646_ (.VDD(vdd),
    .VSS(vss),
    .A(_0048_),
    .B(_0086_),
    .Y(_0087_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0647_ (.VDD(vdd),
    .VSS(vss),
    .A(net15),
    .Y(_0088_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0648_ (.VDD(vdd),
    .VSS(vss),
    .A(_0088_),
    .Y(_0089_));
 gf180mcu_osu_sc_gp9t3v3__aoi22_1 _0649_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0422_),
    .A1(_0047_),
    .B0(_0089_),
    .B1(_0413_),
    .Y(_0090_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0650_ (.VDD(vdd),
    .VSS(vss),
    .A(_0087_),
    .B(_0090_),
    .Y(_0091_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0651_ (.VDD(vdd),
    .VSS(vss),
    .A(_0085_),
    .B(_0091_),
    .Y(_0092_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0652_ (.VDD(vdd),
    .VSS(vss),
    .A(net6),
    .Y(_0093_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0653_ (.VDD(vdd),
    .VSS(vss),
    .A(net10),
    .B(_0093_),
    .Y(_0094_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0654_ (.VDD(vdd),
    .VSS(vss),
    .A(net9),
    .B(net7),
    .Y(_0095_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0655_ (.VDD(vdd),
    .VSS(vss),
    .A(net29),
    .B(_0095_),
    .Y(_0096_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0656_ (.VDD(vdd),
    .VSS(vss),
    .A(_0094_),
    .B(_0096_),
    .Y(_0097_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0657_ (.VDD(vdd),
    .VSS(vss),
    .A(net28),
    .B(_0054_),
    .Y(_0098_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0658_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0053_),
    .A1(_0055_),
    .B(_0098_),
    .Y(_0099_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0659_ (.VDD(vdd),
    .VSS(vss),
    .A(_0097_),
    .B(_0099_),
    .Y(_0100_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0660_ (.VDD(vdd),
    .VSS(vss),
    .A(_0451_),
    .B(_0060_),
    .Y(_0101_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0661_ (.VDD(vdd),
    .VSS(vss),
    .A(_0063_),
    .B(_0052_),
    .Y(_0102_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0662_ (.VDD(vdd),
    .VSS(vss),
    .A(_0082_),
    .B(_0102_),
    .Y(_0103_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0663_ (.VDD(vdd),
    .VSS(vss),
    .A(_0101_),
    .B(_0103_),
    .Y(_0104_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0664_ (.VDD(vdd),
    .VSS(vss),
    .A(_0100_),
    .B(_0104_),
    .Y(_0105_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0665_ (.VDD(vdd),
    .VSS(vss),
    .A(_0056_),
    .B(_0058_),
    .Y(_0106_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0666_ (.VDD(vdd),
    .VSS(vss),
    .A(_0066_),
    .Y(_0107_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0667_ (.VDD(vdd),
    .VSS(vss),
    .A(_0056_),
    .B(_0058_),
    .Y(_0108_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0668_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0106_),
    .A1(_0107_),
    .B(_0108_),
    .Y(_0109_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0669_ (.VDD(vdd),
    .VSS(vss),
    .A(_0105_),
    .B(_0109_),
    .Y(_0110_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0670_ (.VDD(vdd),
    .VSS(vss),
    .A(_0092_),
    .B(_0110_),
    .Y(_0111_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0671_ (.VDD(vdd),
    .VSS(vss),
    .A(_0067_),
    .B(_0069_),
    .Y(_0112_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0672_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0051_),
    .A1(_0070_),
    .B(_0112_),
    .Y(_0113_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0673_ (.VDD(vdd),
    .VSS(vss),
    .A(_0111_),
    .B(_0113_),
    .Y(_0114_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0674_ (.VDD(vdd),
    .VSS(vss),
    .A(_0050_),
    .B(_0114_),
    .Y(_0115_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0675_ (.VDD(vdd),
    .VSS(vss),
    .A(_0080_),
    .B(_0115_),
    .Y(_0116_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0676_ (.VDD(vdd),
    .VSS(vss),
    .A(_0042_),
    .B(_0074_),
    .Y(_0117_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0677_ (.VDD(vdd),
    .VSS(vss),
    .A(_0075_),
    .B(_0077_),
    .Y(_0118_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0678_ (.VDD(vdd),
    .VSS(vss),
    .A(_0117_),
    .B(_0118_),
    .Y(_0119_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0679_ (.VDD(vdd),
    .VSS(vss),
    .A(_0116_),
    .B(_0119_),
    .Y(_0120_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0680_ (.VDD(vdd),
    .VSS(vss),
    .A(_0120_),
    .Y(_0012_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0681_ (.VDD(vdd),
    .VSS(vss),
    .A(_0111_),
    .B(_0113_),
    .Y(_0121_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0682_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0050_),
    .A1(_0114_),
    .B(_0121_),
    .Y(_0122_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0683_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0083_),
    .A1(_0084_),
    .B(_0091_),
    .Y(_0123_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0684_ (.VDD(vdd),
    .VSS(vss),
    .A(_0081_),
    .B(_0052_),
    .Y(_0124_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0685_ (.VDD(vdd),
    .VSS(vss),
    .A(_0064_),
    .B(_0124_),
    .Y(_0125_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0686_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0101_),
    .A1(_0103_),
    .B(_0125_),
    .Y(_0126_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0687_ (.VDD(vdd),
    .VSS(vss),
    .A(net16),
    .Y(_0127_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0688_ (.VDD(vdd),
    .VSS(vss),
    .A(_0412_),
    .B(_0127_),
    .Y(_0128_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0689_ (.VDD(vdd),
    .VSS(vss),
    .A(_0433_),
    .B(_0046_),
    .Y(_0129_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0690_ (.VDD(vdd),
    .VSS(vss),
    .A(_0086_),
    .B(_0129_),
    .Y(_0130_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0691_ (.VDD(vdd),
    .VSS(vss),
    .A(_0128_),
    .B(_0130_),
    .Y(_0131_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0692_ (.VDD(vdd),
    .VSS(vss),
    .A(_0126_),
    .B(_0131_),
    .Y(_0132_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0693_ (.VDD(vdd),
    .VSS(vss),
    .A(_0087_),
    .B(_0132_),
    .Y(_0133_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0694_ (.VDD(vdd),
    .VSS(vss),
    .A(net4),
    .Y(_0134_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0695_ (.VDD(vdd),
    .VSS(vss),
    .A(_0134_),
    .B(_0034_),
    .Y(_0135_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0696_ (.VDD(vdd),
    .VSS(vss),
    .A(_0093_),
    .Y(_0136_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0697_ (.VDD(vdd),
    .VSS(vss),
    .A(_0063_),
    .B(_0136_),
    .Y(_0137_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0698_ (.VDD(vdd),
    .VSS(vss),
    .A(_0124_),
    .B(_0137_),
    .Y(_0138_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0699_ (.VDD(vdd),
    .VSS(vss),
    .A(_0135_),
    .B(_0138_),
    .Y(_0139_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0700_ (.VDD(vdd),
    .VSS(vss),
    .A(net7),
    .Y(_0140_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0701_ (.VDD(vdd),
    .VSS(vss),
    .A(_0419_),
    .B(_0140_),
    .Y(_0141_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0702_ (.VDD(vdd),
    .VSS(vss),
    .A(_0405_),
    .B(net8),
    .Y(_0142_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0703_ (.VDD(vdd),
    .VSS(vss),
    .A(net30),
    .B(_0142_),
    .Y(_0143_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0704_ (.VDD(vdd),
    .VSS(vss),
    .A(_0141_),
    .B(_0143_),
    .Y(_0144_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0705_ (.VDD(vdd),
    .VSS(vss),
    .A(net29),
    .B(_0095_),
    .Y(_0145_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0706_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0094_),
    .A1(_0096_),
    .B(_0145_),
    .Y(_0146_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0707_ (.VDD(vdd),
    .VSS(vss),
    .A(_0144_),
    .B(_0146_),
    .Y(_0147_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0708_ (.VDD(vdd),
    .VSS(vss),
    .A(_0139_),
    .B(_0147_),
    .Y(_0148_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0709_ (.VDD(vdd),
    .VSS(vss),
    .A(_0104_),
    .Y(_0149_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0710_ (.VDD(vdd),
    .VSS(vss),
    .A(_0097_),
    .B(_0099_),
    .Y(_0150_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0711_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0100_),
    .A1(_0149_),
    .B(_0150_),
    .Y(_0151_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0712_ (.VDD(vdd),
    .VSS(vss),
    .A(_0148_),
    .B(_0151_),
    .Y(_0152_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0713_ (.VDD(vdd),
    .VSS(vss),
    .A(_0133_),
    .B(_0152_),
    .Y(_0153_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0714_ (.VDD(vdd),
    .VSS(vss),
    .A(_0105_),
    .B(_0109_),
    .Y(_0154_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0715_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0092_),
    .A1(_0110_),
    .B(_0154_),
    .Y(_0155_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0716_ (.VDD(vdd),
    .VSS(vss),
    .A(_0153_),
    .B(_0155_),
    .Y(_0156_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0717_ (.VDD(vdd),
    .VSS(vss),
    .A(_0123_),
    .B(_0156_),
    .Y(_0157_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0718_ (.VDD(vdd),
    .VSS(vss),
    .A(_0122_),
    .B(_0157_),
    .Y(_0158_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0719_ (.VDD(vdd),
    .VSS(vss),
    .A(_0122_),
    .B(_0157_),
    .Y(_0159_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0720_ (.VDD(vdd),
    .VSS(vss),
    .A(_0158_),
    .B(_0159_),
    .Y(_0160_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0721_ (.VDD(vdd),
    .VSS(vss),
    .A(_0080_),
    .B(_0115_),
    .Y(_0161_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0722_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0117_),
    .A1(_0118_),
    .B(_0116_),
    .Y(_0162_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0723_ (.VDD(vdd),
    .VSS(vss),
    .A(_0161_),
    .B(_0162_),
    .Y(_0163_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0724_ (.VDD(vdd),
    .VSS(vss),
    .A(_0160_),
    .B(_0163_),
    .Y(_0164_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0725_ (.VDD(vdd),
    .VSS(vss),
    .A(_0164_),
    .Y(_0013_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0726_ (.VDD(vdd),
    .VSS(vss),
    .A(_0153_),
    .B(_0155_),
    .Y(_0165_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0727_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0123_),
    .A1(_0156_),
    .B(_0165_),
    .Y(_0166_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0728_ (.VDD(vdd),
    .VSS(vss),
    .A(_0131_),
    .Y(_0167_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0729_ (.VDD(vdd),
    .VSS(vss),
    .A(_0126_),
    .B(_0167_),
    .Y(_0168_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0730_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0087_),
    .A1(_0132_),
    .B(_0168_),
    .Y(_0169_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0731_ (.VDD(vdd),
    .VSS(vss),
    .A(_0148_),
    .B(_0151_),
    .Y(_0170_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0732_ (.VDD(vdd),
    .VSS(vss),
    .A(_0148_),
    .B(_0151_),
    .Y(_0171_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0733_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0133_),
    .A1(_0170_),
    .B(_0171_),
    .Y(_0172_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0734_ (.VDD(vdd),
    .VSS(vss),
    .A(_0086_),
    .B(_0129_),
    .Y(_0173_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0735_ (.VDD(vdd),
    .VSS(vss),
    .A(_0128_),
    .B(_0130_),
    .Y(_0174_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0736_ (.VDD(vdd),
    .VSS(vss),
    .A(_0173_),
    .B(_0174_),
    .Y(_0175_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0737_ (.VDD(vdd),
    .VSS(vss),
    .A(_0175_),
    .Y(_0176_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0738_ (.VDD(vdd),
    .VSS(vss),
    .A(_0081_),
    .B(_0093_),
    .Y(_0177_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0739_ (.VDD(vdd),
    .VSS(vss),
    .A(_0102_),
    .B(_0177_),
    .Y(_0178_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0740_ (.VDD(vdd),
    .VSS(vss),
    .A(_0135_),
    .B(_0138_),
    .Y(_0179_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0741_ (.VDD(vdd),
    .VSS(vss),
    .A(_0178_),
    .B(_0179_),
    .Y(_0180_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0742_ (.VDD(vdd),
    .VSS(vss),
    .A(net16),
    .Y(_0181_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0743_ (.VDD(vdd),
    .VSS(vss),
    .A(_0422_),
    .B(_0181_),
    .Y(_0182_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0744_ (.VDD(vdd),
    .VSS(vss),
    .A(_0134_),
    .B(_0088_),
    .Y(_0183_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0745_ (.VDD(vdd),
    .VSS(vss),
    .A(_0129_),
    .B(_0183_),
    .Y(_0184_));
 gf180mcu_osu_sc_gp9t3v3__aoi22_1 _0746_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0134_),
    .A1(_0047_),
    .B0(_0089_),
    .B1(_0451_),
    .Y(_0185_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0747_ (.VDD(vdd),
    .VSS(vss),
    .A(_0184_),
    .B(_0185_),
    .Y(_0186_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0748_ (.VDD(vdd),
    .VSS(vss),
    .A(_0182_),
    .B(_0186_),
    .Y(_0187_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0749_ (.VDD(vdd),
    .VSS(vss),
    .A(_0180_),
    .B(_0187_),
    .Y(_0188_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0750_ (.VDD(vdd),
    .VSS(vss),
    .A(_0176_),
    .B(_0188_),
    .Y(_0189_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0751_ (.VDD(vdd),
    .VSS(vss),
    .A(_0139_),
    .Y(_0190_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0752_ (.VDD(vdd),
    .VSS(vss),
    .A(_0144_),
    .B(_0146_),
    .Y(_0191_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0753_ (.VDD(vdd),
    .VSS(vss),
    .A(_0144_),
    .B(_0146_),
    .Y(_0192_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0754_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0190_),
    .A1(_0191_),
    .B(_0192_),
    .Y(_0193_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0755_ (.VDD(vdd),
    .VSS(vss),
    .A(_0052_),
    .Y(_0194_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0756_ (.VDD(vdd),
    .VSS(vss),
    .A(_0194_),
    .B(_0060_),
    .Y(_0195_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0757_ (.VDD(vdd),
    .VSS(vss),
    .A(_0430_),
    .B(_0140_),
    .Y(_0196_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0758_ (.VDD(vdd),
    .VSS(vss),
    .A(_0177_),
    .B(_0196_),
    .Y(_0197_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0759_ (.VDD(vdd),
    .VSS(vss),
    .A(_0195_),
    .B(_0197_),
    .Y(_0198_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0760_ (.VDD(vdd),
    .VSS(vss),
    .A(net31),
    .Y(_0199_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0761_ (.VDD(vdd),
    .VSS(vss),
    .A(net8),
    .Y(_0200_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0762_ (.VDD(vdd),
    .VSS(vss),
    .A(_0418_),
    .B(_0200_),
    .Y(_0201_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0763_ (.VDD(vdd),
    .VSS(vss),
    .A(_0199_),
    .B(_0201_),
    .Y(_0202_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0764_ (.VDD(vdd),
    .VSS(vss),
    .A(_0202_),
    .Y(_0203_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0765_ (.VDD(vdd),
    .VSS(vss),
    .A(net30),
    .B(_0142_),
    .Y(_0204_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0766_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0141_),
    .A1(_0143_),
    .B(_0204_),
    .Y(_0205_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0767_ (.VDD(vdd),
    .VSS(vss),
    .A(_0203_),
    .B(_0205_),
    .Y(_0206_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0768_ (.VDD(vdd),
    .VSS(vss),
    .A(_0198_),
    .B(_0206_),
    .Y(_0207_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0769_ (.VDD(vdd),
    .VSS(vss),
    .A(_0193_),
    .B(_0207_),
    .Y(_0208_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0770_ (.VDD(vdd),
    .VSS(vss),
    .A(_0189_),
    .B(_0208_),
    .Y(_0209_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0771_ (.VDD(vdd),
    .VSS(vss),
    .A(_0172_),
    .B(_0209_),
    .Y(_0210_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0772_ (.VDD(vdd),
    .VSS(vss),
    .A(_0169_),
    .B(_0210_),
    .Y(_0211_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0773_ (.VDD(vdd),
    .VSS(vss),
    .A(_0166_),
    .B(_0211_),
    .Y(_0212_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0774_ (.VDD(vdd),
    .VSS(vss),
    .A(_0158_),
    .Y(_0213_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0775_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0213_),
    .A1(_0163_),
    .B(_0159_),
    .Y(_0214_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0776_ (.VDD(vdd),
    .VSS(vss),
    .A(_0212_),
    .B(_0214_),
    .Y(_0215_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0777_ (.VDD(vdd),
    .VSS(vss),
    .A(_0215_),
    .Y(_0014_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0778_ (.VDD(vdd),
    .VSS(vss),
    .A(_0172_),
    .B(_0209_),
    .Y(_0216_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0779_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0169_),
    .A1(_0210_),
    .B(_0216_),
    .Y(_0217_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0780_ (.VDD(vdd),
    .VSS(vss),
    .A(_0187_),
    .Y(_0218_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0781_ (.VDD(vdd),
    .VSS(vss),
    .A(_0180_),
    .B(_0218_),
    .Y(_0219_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0782_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0176_),
    .A1(_0188_),
    .B(_0219_),
    .Y(_0220_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0783_ (.VDD(vdd),
    .VSS(vss),
    .A(_0193_),
    .B(_0207_),
    .Y(_0221_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0784_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0189_),
    .A1(_0208_),
    .B(_0221_),
    .Y(_0222_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0785_ (.VDD(vdd),
    .VSS(vss),
    .A(_0182_),
    .B(_0186_),
    .Y(_0223_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0786_ (.VDD(vdd),
    .VSS(vss),
    .A(_0184_),
    .B(_0223_),
    .Y(_0224_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0787_ (.VDD(vdd),
    .VSS(vss),
    .A(_0081_),
    .B(net7),
    .Y(_0225_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0788_ (.VDD(vdd),
    .VSS(vss),
    .A(_0225_),
    .Y(_0226_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0789_ (.VDD(vdd),
    .VSS(vss),
    .A(_0137_),
    .B(_0226_),
    .Y(_0227_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0790_ (.VDD(vdd),
    .VSS(vss),
    .A(_0195_),
    .B(_0197_),
    .Y(_0228_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0791_ (.VDD(vdd),
    .VSS(vss),
    .A(_0227_),
    .B(_0228_),
    .Y(_0229_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0792_ (.VDD(vdd),
    .VSS(vss),
    .A(_0451_),
    .B(_0127_),
    .Y(_0230_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0793_ (.VDD(vdd),
    .VSS(vss),
    .A(_0194_),
    .B(_0046_),
    .Y(_0231_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0794_ (.VDD(vdd),
    .VSS(vss),
    .A(_0183_),
    .B(_0231_),
    .Y(_0232_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0795_ (.VDD(vdd),
    .VSS(vss),
    .A(_0230_),
    .B(_0232_),
    .Y(_0233_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0796_ (.VDD(vdd),
    .VSS(vss),
    .A(_0229_),
    .B(_0233_),
    .Y(_0234_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0797_ (.VDD(vdd),
    .VSS(vss),
    .A(_0224_),
    .B(_0234_),
    .Y(_0235_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0798_ (.VDD(vdd),
    .VSS(vss),
    .A(_0203_),
    .B(_0205_),
    .Y(_0236_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0799_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0198_),
    .A1(_0206_),
    .B(_0236_),
    .Y(_0237_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0800_ (.VDD(vdd),
    .VSS(vss),
    .A(_0136_),
    .B(net13),
    .Y(_0238_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0801_ (.VDD(vdd),
    .VSS(vss),
    .A(_0063_),
    .B(net8),
    .Y(_0239_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0802_ (.VDD(vdd),
    .VSS(vss),
    .A(_0225_),
    .B(_0239_),
    .Y(_0240_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0803_ (.VDD(vdd),
    .VSS(vss),
    .A(_0238_),
    .B(_0240_),
    .Y(_0241_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0804_ (.VDD(vdd),
    .VSS(vss),
    .A(_0199_),
    .B(_0201_),
    .Y(_0242_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0805_ (.VDD(vdd),
    .VSS(vss),
    .A(net32),
    .B(_0242_),
    .Y(_0243_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0806_ (.VDD(vdd),
    .VSS(vss),
    .A(_0241_),
    .B(_0243_),
    .Y(_0244_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0807_ (.VDD(vdd),
    .VSS(vss),
    .A(_0244_),
    .Y(_0245_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0808_ (.VDD(vdd),
    .VSS(vss),
    .A(_0237_),
    .B(_0245_),
    .Y(_0246_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0809_ (.VDD(vdd),
    .VSS(vss),
    .A(_0235_),
    .B(_0246_),
    .Y(_0247_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0810_ (.VDD(vdd),
    .VSS(vss),
    .A(_0222_),
    .B(_0247_),
    .Y(_0248_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0811_ (.VDD(vdd),
    .VSS(vss),
    .A(_0220_),
    .B(_0248_),
    .Y(_0249_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0812_ (.VDD(vdd),
    .VSS(vss),
    .A(_0217_),
    .B(_0249_),
    .Y(_0250_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0813_ (.VDD(vdd),
    .VSS(vss),
    .A(_0159_),
    .Y(_0251_));
 gf180mcu_osu_sc_gp9t3v3__oai31_1 _0814_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0161_),
    .A1(_0162_),
    .A2(_0251_),
    .B(_0158_),
    .Y(_0252_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0815_ (.VDD(vdd),
    .VSS(vss),
    .A(_0166_),
    .B(_0211_),
    .Y(_0253_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0816_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0212_),
    .A1(_0252_),
    .B(_0253_),
    .Y(_0254_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0817_ (.VDD(vdd),
    .VSS(vss),
    .A(_0250_),
    .B(_0254_),
    .Y(_0255_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0818_ (.VDD(vdd),
    .VSS(vss),
    .A(_0255_),
    .Y(_0015_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0819_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0227_),
    .A1(_0228_),
    .B(_0233_),
    .Y(_0256_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0820_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0184_),
    .A1(_0223_),
    .B(_0234_),
    .Y(_0257_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0821_ (.VDD(vdd),
    .VSS(vss),
    .A(_0256_),
    .B(_0257_),
    .Y(_0258_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0822_ (.VDD(vdd),
    .VSS(vss),
    .A(_0183_),
    .B(_0231_),
    .Y(_0259_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0823_ (.VDD(vdd),
    .VSS(vss),
    .A(_0230_),
    .B(_0232_),
    .Y(_0260_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0824_ (.VDD(vdd),
    .VSS(vss),
    .A(_0259_),
    .B(_0260_),
    .Y(_0261_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0825_ (.VDD(vdd),
    .VSS(vss),
    .A(_0238_),
    .Y(_0262_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0826_ (.VDD(vdd),
    .VSS(vss),
    .A(_0226_),
    .B(_0239_),
    .Y(_0263_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0827_ (.VDD(vdd),
    .VSS(vss),
    .A(_0226_),
    .B(_0239_),
    .Y(_0264_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0828_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0262_),
    .A1(_0263_),
    .B(_0264_),
    .Y(_0265_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0829_ (.VDD(vdd),
    .VSS(vss),
    .A(_0134_),
    .B(_0127_),
    .Y(_0266_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0830_ (.VDD(vdd),
    .VSS(vss),
    .A(_0194_),
    .B(_0088_),
    .Y(_0267_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0831_ (.VDD(vdd),
    .VSS(vss),
    .A(_0093_),
    .B(net14),
    .Y(_0268_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0832_ (.VDD(vdd),
    .VSS(vss),
    .A(_0267_),
    .B(_0268_),
    .Y(_0269_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0833_ (.VDD(vdd),
    .VSS(vss),
    .A(_0266_),
    .B(_0269_),
    .Y(_0270_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0834_ (.VDD(vdd),
    .VSS(vss),
    .A(_0265_),
    .B(_0270_),
    .Y(_0271_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0835_ (.VDD(vdd),
    .VSS(vss),
    .A(_0261_),
    .B(_0271_),
    .Y(_0272_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0836_ (.VDD(vdd),
    .VSS(vss),
    .A(_0060_),
    .B(_0200_),
    .Y(_0273_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0837_ (.VDD(vdd),
    .VSS(vss),
    .A(_0226_),
    .B(_0273_),
    .Y(_0274_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0838_ (.VDD(vdd),
    .VSS(vss),
    .A(_0140_),
    .Y(_0275_));
 gf180mcu_osu_sc_gp9t3v3__aoi22_1 _0839_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0034_),
    .A1(_0275_),
    .B0(_0200_),
    .B1(_0446_),
    .Y(_0276_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0840_ (.VDD(vdd),
    .VSS(vss),
    .A(_0274_),
    .B(_0276_),
    .Y(_0277_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0841_ (.VDD(vdd),
    .VSS(vss),
    .A(net18),
    .B(_0277_),
    .Y(_0278_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0842_ (.VDD(vdd),
    .VSS(vss),
    .A(net32),
    .B(_0242_),
    .Y(_0279_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0843_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0241_),
    .A1(_0243_),
    .B(_0279_),
    .Y(_0280_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0844_ (.VDD(vdd),
    .VSS(vss),
    .A(_0278_),
    .B(_0280_),
    .Y(_0281_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0845_ (.VDD(vdd),
    .VSS(vss),
    .A(_0272_),
    .B(_0281_),
    .Y(_0282_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0846_ (.VDD(vdd),
    .VSS(vss),
    .A(_0237_),
    .B(_0245_),
    .Y(_0283_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0847_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0235_),
    .A1(_0246_),
    .B(_0283_),
    .Y(_0284_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0848_ (.VDD(vdd),
    .VSS(vss),
    .A(_0282_),
    .B(_0284_),
    .Y(_0285_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0849_ (.VDD(vdd),
    .VSS(vss),
    .A(_0258_),
    .B(_0285_),
    .Y(_0286_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0850_ (.VDD(vdd),
    .VSS(vss),
    .A(_0220_),
    .Y(_0287_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0851_ (.VDD(vdd),
    .VSS(vss),
    .A(_0189_),
    .B(_0208_),
    .Y(_0288_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0852_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0221_),
    .A1(_0288_),
    .B(_0247_),
    .Y(_0289_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0853_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0287_),
    .A1(_0248_),
    .B(_0289_),
    .Y(_0290_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0854_ (.VDD(vdd),
    .VSS(vss),
    .A(_0286_),
    .B(_0290_),
    .Y(_0291_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0855_ (.VDD(vdd),
    .VSS(vss),
    .A(_0212_),
    .B(_0250_),
    .Y(_0292_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0856_ (.VDD(vdd),
    .VSS(vss),
    .A(_0217_),
    .B(_0249_),
    .Y(_0293_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0857_ (.VDD(vdd),
    .VSS(vss),
    .A(_0217_),
    .B(_0249_),
    .Y(_0294_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0858_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0253_),
    .A1(_0293_),
    .B(_0294_),
    .Y(_0295_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0859_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0214_),
    .A1(_0292_),
    .B(_0295_),
    .Y(_0296_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0860_ (.VDD(vdd),
    .VSS(vss),
    .A(_0291_),
    .B(_0296_),
    .Y(_0297_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0861_ (.VDD(vdd),
    .VSS(vss),
    .A(_0297_),
    .Y(_0005_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0862_ (.VDD(vdd),
    .VSS(vss),
    .A(_0265_),
    .Y(_0298_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0863_ (.VDD(vdd),
    .VSS(vss),
    .A(_0298_),
    .B(_0270_),
    .Y(_0299_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0864_ (.VDD(vdd),
    .VSS(vss),
    .A(_0298_),
    .B(_0270_),
    .Y(_0300_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0865_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0261_),
    .A1(_0299_),
    .B(_0300_),
    .Y(_0301_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0866_ (.VDD(vdd),
    .VSS(vss),
    .A(net18),
    .B(_0277_),
    .Y(_0302_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0867_ (.VDD(vdd),
    .VSS(vss),
    .A(_0200_),
    .Y(_0303_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0868_ (.VDD(vdd),
    .VSS(vss),
    .A(_0034_),
    .B(_0303_),
    .Y(_0304_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0869_ (.VDD(vdd),
    .VSS(vss),
    .A(net19),
    .B(_0304_),
    .Y(_0305_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0870_ (.VDD(vdd),
    .VSS(vss),
    .A(_0302_),
    .B(_0305_),
    .Y(_0306_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0871_ (.VDD(vdd),
    .VSS(vss),
    .A(_0267_),
    .B(_0268_),
    .Y(_0307_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0872_ (.VDD(vdd),
    .VSS(vss),
    .A(_0266_),
    .B(_0269_),
    .Y(_0308_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0873_ (.VDD(vdd),
    .VSS(vss),
    .A(_0307_),
    .B(_0308_),
    .Y(_0309_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0874_ (.VDD(vdd),
    .VSS(vss),
    .A(_0194_),
    .B(_0127_),
    .Y(_0310_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0875_ (.VDD(vdd),
    .VSS(vss),
    .A(_0140_),
    .B(net15),
    .Y(_0311_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0876_ (.VDD(vdd),
    .VSS(vss),
    .A(_0268_),
    .B(_0311_),
    .Y(_0312_));
 gf180mcu_osu_sc_gp9t3v3__aoi22_1 _0877_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0046_),
    .A1(_0275_),
    .B0(_0088_),
    .B1(_0136_),
    .Y(_0313_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0878_ (.VDD(vdd),
    .VSS(vss),
    .A(_0312_),
    .B(_0313_),
    .Y(_0314_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0879_ (.VDD(vdd),
    .VSS(vss),
    .A(_0310_),
    .B(_0314_),
    .Y(_0315_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0880_ (.VDD(vdd),
    .VSS(vss),
    .A(_0274_),
    .B(_0315_),
    .Y(_0316_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0881_ (.VDD(vdd),
    .VSS(vss),
    .A(_0309_),
    .B(_0316_),
    .Y(_0317_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0882_ (.VDD(vdd),
    .VSS(vss),
    .A(_0306_),
    .B(_0317_),
    .Y(_0318_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0883_ (.VDD(vdd),
    .VSS(vss),
    .A(_0241_),
    .B(_0243_),
    .Y(_0319_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0884_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0279_),
    .A1(_0319_),
    .B(_0278_),
    .Y(_0320_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0885_ (.VDD(vdd),
    .VSS(vss),
    .A(_0272_),
    .B(_0281_),
    .Y(_0321_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0886_ (.VDD(vdd),
    .VSS(vss),
    .A(_0320_),
    .B(_0321_),
    .Y(_0322_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0887_ (.VDD(vdd),
    .VSS(vss),
    .A(_0318_),
    .B(_0322_),
    .Y(_0323_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0888_ (.VDD(vdd),
    .VSS(vss),
    .A(_0301_),
    .B(_0323_),
    .Y(_0324_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0889_ (.VDD(vdd),
    .VSS(vss),
    .A(_0282_),
    .B(_0284_),
    .Y(_0325_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0890_ (.VDD(vdd),
    .VSS(vss),
    .A(_0282_),
    .B(_0284_),
    .Y(_0326_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0891_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0258_),
    .A1(_0325_),
    .B(_0326_),
    .Y(_0327_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0892_ (.VDD(vdd),
    .VSS(vss),
    .A(_0324_),
    .B(_0327_),
    .Y(_0328_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0893_ (.VDD(vdd),
    .VSS(vss),
    .A(_0286_),
    .B(_0290_),
    .Y(_0329_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0894_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0291_),
    .A1(_0296_),
    .B(_0329_),
    .Y(_0330_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0895_ (.VDD(vdd),
    .VSS(vss),
    .A(_0328_),
    .B(_0330_),
    .Y(_0331_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0896_ (.VDD(vdd),
    .VSS(vss),
    .A(_0331_),
    .Y(_0006_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0897_ (.VDD(vdd),
    .VSS(vss),
    .A(_0274_),
    .B(_0315_),
    .Y(_0332_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0898_ (.VDD(vdd),
    .VSS(vss),
    .A(_0274_),
    .B(_0315_),
    .Y(_0333_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0899_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0309_),
    .A1(_0332_),
    .B(_0333_),
    .Y(_0334_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0900_ (.VDD(vdd),
    .VSS(vss),
    .A(_0306_),
    .B(_0317_),
    .Y(_0335_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0901_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0302_),
    .A1(_0305_),
    .B(_0335_),
    .Y(_0336_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0902_ (.VDD(vdd),
    .VSS(vss),
    .A(net19),
    .B(_0304_),
    .Y(_0337_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0903_ (.VDD(vdd),
    .VSS(vss),
    .A(net20),
    .B(_0337_),
    .Y(_0338_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0904_ (.VDD(vdd),
    .VSS(vss),
    .A(_0136_),
    .B(_0181_),
    .Y(_0339_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0905_ (.VDD(vdd),
    .VSS(vss),
    .A(_0047_),
    .B(_0303_),
    .Y(_0340_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0906_ (.VDD(vdd),
    .VSS(vss),
    .A(_0311_),
    .B(_0340_),
    .Y(_0341_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0907_ (.VDD(vdd),
    .VSS(vss),
    .A(_0339_),
    .B(_0341_),
    .Y(_0342_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0908_ (.VDD(vdd),
    .VSS(vss),
    .A(_0310_),
    .B(_0314_),
    .Y(_0343_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0909_ (.VDD(vdd),
    .VSS(vss),
    .A(_0312_),
    .B(_0343_),
    .Y(_0344_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0910_ (.VDD(vdd),
    .VSS(vss),
    .A(_0342_),
    .B(_0344_),
    .Y(_0345_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0911_ (.VDD(vdd),
    .VSS(vss),
    .A(_0338_),
    .B(_0345_),
    .Y(_0346_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0912_ (.VDD(vdd),
    .VSS(vss),
    .A(_0336_),
    .B(_0346_),
    .Y(_0347_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0913_ (.VDD(vdd),
    .VSS(vss),
    .A(_0334_),
    .B(_0347_),
    .Y(_0348_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0914_ (.VDD(vdd),
    .VSS(vss),
    .A(_0318_),
    .B(_0322_),
    .Y(_0349_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0915_ (.VDD(vdd),
    .VSS(vss),
    .A(_0318_),
    .B(_0322_),
    .Y(_0350_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0916_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0301_),
    .A1(_0349_),
    .B(_0350_),
    .Y(_0351_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0917_ (.VDD(vdd),
    .VSS(vss),
    .A(_0348_),
    .B(_0351_),
    .Y(_0352_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0918_ (.VDD(vdd),
    .VSS(vss),
    .A(_0292_),
    .Y(_0353_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0919_ (.VDD(vdd),
    .VSS(vss),
    .A(_0291_),
    .B(_0328_),
    .Y(_0354_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0920_ (.VDD(vdd),
    .VSS(vss),
    .A(_0324_),
    .B(_0327_),
    .Y(_0355_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0921_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0324_),
    .A1(_0327_),
    .B(_0329_),
    .Y(_0356_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0922_ (.VDD(vdd),
    .VSS(vss),
    .A(_0291_),
    .B(_0328_),
    .Y(_0357_));
 gf180mcu_osu_sc_gp9t3v3__aoi22_1 _0923_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0355_),
    .A1(_0356_),
    .B0(_0357_),
    .B1(_0295_),
    .Y(_0358_));
 gf180mcu_osu_sc_gp9t3v3__oai31_1 _0924_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0252_),
    .A1(_0353_),
    .A2(_0354_),
    .B(_0358_),
    .Y(_0359_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0925_ (.VDD(vdd),
    .VSS(vss),
    .A(_0352_),
    .B(_0359_),
    .Y(_0360_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0926_ (.VDD(vdd),
    .VSS(vss),
    .A(_0360_),
    .Y(_0007_));
 gf180mcu_osu_sc_gp9t3v3__oai21_1 _0927_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0312_),
    .A1(_0343_),
    .B(_0342_),
    .Y(_0361_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0928_ (.VDD(vdd),
    .VSS(vss),
    .A(_0311_),
    .B(_0340_),
    .Y(_0362_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0929_ (.VDD(vdd),
    .VSS(vss),
    .A(_0339_),
    .B(_0341_),
    .Y(_0363_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0930_ (.VDD(vdd),
    .VSS(vss),
    .A(_0362_),
    .B(_0363_),
    .Y(_0364_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0931_ (.VDD(vdd),
    .VSS(vss),
    .A(_0089_),
    .B(_0303_),
    .Y(_0365_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0932_ (.VDD(vdd),
    .VSS(vss),
    .A(_0275_),
    .B(_0181_),
    .Y(_0366_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0933_ (.VDD(vdd),
    .VSS(vss),
    .A(_0365_),
    .B(_0366_),
    .Y(_0367_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0934_ (.VDD(vdd),
    .VSS(vss),
    .A(_0364_),
    .B(_0367_),
    .Y(_0368_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0935_ (.VDD(vdd),
    .VSS(vss),
    .A(net21),
    .B(_0368_),
    .Y(_0369_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0936_ (.VDD(vdd),
    .VSS(vss),
    .A(net20),
    .B(_0337_),
    .Y(_0370_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0937_ (.VDD(vdd),
    .VSS(vss),
    .A(_0338_),
    .Y(_0371_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0938_ (.VDD(vdd),
    .VSS(vss),
    .A(_0371_),
    .B(_0345_),
    .Y(_0372_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0939_ (.VDD(vdd),
    .VSS(vss),
    .A(_0370_),
    .B(_0372_),
    .Y(_0373_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0940_ (.VDD(vdd),
    .VSS(vss),
    .A(_0369_),
    .B(_0373_),
    .Y(_0374_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0941_ (.VDD(vdd),
    .VSS(vss),
    .A(_0361_),
    .B(_0374_),
    .Y(_0375_));
 gf180mcu_osu_sc_gp9t3v3__and2_1 _0942_ (.VDD(vdd),
    .VSS(vss),
    .A(_0334_),
    .B(_0347_),
    .Y(_0376_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0943_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0336_),
    .A1(_0346_),
    .B(_0376_),
    .Y(_0377_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0944_ (.VDD(vdd),
    .VSS(vss),
    .A(_0375_),
    .B(_0377_),
    .Y(_0378_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0945_ (.VDD(vdd),
    .VSS(vss),
    .A(_0378_),
    .Y(_0379_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0946_ (.VDD(vdd),
    .VSS(vss),
    .A(_0375_),
    .B(_0377_),
    .Y(_0380_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0947_ (.VDD(vdd),
    .VSS(vss),
    .A(_0379_),
    .B(_0380_),
    .Y(_0381_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0948_ (.VDD(vdd),
    .VSS(vss),
    .A(_0348_),
    .B(_0351_),
    .Y(_0382_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0949_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0352_),
    .A1(_0359_),
    .B(_0382_),
    .Y(_0383_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0950_ (.VDD(vdd),
    .VSS(vss),
    .A(_0381_),
    .B(_0383_),
    .Y(_0384_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0951_ (.VDD(vdd),
    .VSS(vss),
    .A(_0384_),
    .Y(_0008_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0952_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0370_),
    .A1(_0372_),
    .B(_0369_),
    .Y(_0385_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0953_ (.VDD(vdd),
    .VSS(vss),
    .A(_0361_),
    .B(_0374_),
    .Y(_0386_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0954_ (.VDD(vdd),
    .VSS(vss),
    .A(_0385_),
    .B(_0386_),
    .Y(_0387_));
 gf180mcu_osu_sc_gp9t3v3__or2_1 _0955_ (.VDD(vdd),
    .VSS(vss),
    .A(_0364_),
    .B(_0367_),
    .Y(_0388_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0956_ (.VDD(vdd),
    .VSS(vss),
    .A(net21),
    .B(_0368_),
    .Y(_0389_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0957_ (.VDD(vdd),
    .VSS(vss),
    .A(_0388_),
    .B(_0389_),
    .Y(_0390_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0958_ (.VDD(vdd),
    .VSS(vss),
    .A(_0303_),
    .B(_0181_),
    .Y(_0391_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0959_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0275_),
    .A1(_0089_),
    .B(_0391_),
    .Y(_0392_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0960_ (.VDD(vdd),
    .VSS(vss),
    .A(net22),
    .B(_0392_),
    .Y(_0393_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0961_ (.VDD(vdd),
    .VSS(vss),
    .A(_0390_),
    .B(_0393_),
    .Y(_0394_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0962_ (.VDD(vdd),
    .VSS(vss),
    .A(_0387_),
    .B(_0394_),
    .Y(_0395_));
 gf180mcu_osu_sc_gp9t3v3__nand2_1 _0963_ (.VDD(vdd),
    .VSS(vss),
    .A(_0352_),
    .B(_0359_),
    .Y(_0396_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0964_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0382_),
    .A1(_0378_),
    .B(_0380_),
    .Y(_0397_));
 gf180mcu_osu_sc_gp9t3v3__oai31_1 _0965_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0396_),
    .A1(_0379_),
    .A2(_0380_),
    .B(_0397_),
    .Y(_0398_));
 gf180mcu_osu_sc_gp9t3v3__xor2_1 _0966_ (.VDD(vdd),
    .VSS(vss),
    .A(_0395_),
    .B(_0398_),
    .Y(_0399_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0967_ (.VDD(vdd),
    .VSS(vss),
    .A(_0399_),
    .Y(_0009_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0968_ (.VDD(vdd),
    .VSS(vss),
    .A(_0387_),
    .B(_0394_),
    .Y(_0400_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0969_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0395_),
    .A1(_0398_),
    .B(_0400_),
    .Y(_0401_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0970_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0388_),
    .A1(_0389_),
    .B(_0393_),
    .Y(_0402_));
 gf180mcu_osu_sc_gp9t3v3__clkinv_1 _0971_ (.VDD(vdd),
    .VSS(vss),
    .A(net22),
    .Y(_0403_));
 gf180mcu_osu_sc_gp9t3v3__aoi21_1 _0972_ (.VDD(vdd),
    .VSS(vss),
    .A0(_0403_),
    .A1(_0311_),
    .B(_0391_),
    .Y(_0404_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0973_ (.VDD(vdd),
    .VSS(vss),
    .A(net23),
    .B(_0404_),
    .Y(_0406_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0974_ (.VDD(vdd),
    .VSS(vss),
    .A(_0402_),
    .B(_0406_),
    .Y(_0407_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0975_ (.VDD(vdd),
    .VSS(vss),
    .A(_0401_),
    .B(_0407_),
    .Y(_0408_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0976_ (.VDD(vdd),
    .VSS(vss),
    .A(_0408_),
    .Y(_0010_));
 gf180mcu_osu_sc_gp9t3v3__nor2_1 _0977_ (.VDD(vdd),
    .VSS(vss),
    .A(_0022_),
    .B(_0076_),
    .Y(_0409_));
 gf180mcu_osu_sc_gp9t3v3__xnor2_1 _0978_ (.VDD(vdd),
    .VSS(vss),
    .A(_0041_),
    .B(_0409_),
    .Y(_0410_));
 gf180mcu_osu_sc_gp9t3v3__clkbuf_1 _0979_ (.VDD(vdd),
    .VSS(vss),
    .A(_0410_),
    .Y(_0004_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0980_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net50),
    .D(_0000_),
    .Q(\o_tmp[0][0] ),
    .QN(_0459_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0981_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net51),
    .D(_0001_),
    .Q(\o_tmp[0][1] ),
    .QN(_0460_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0982_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net52),
    .D(_0002_),
    .Q(\o_tmp[0][2] ),
    .QN(_0461_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0983_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net56),
    .D(_0003_),
    .Q(\o_tmp[0][3] ),
    .QN(_0462_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0984_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net57),
    .D(_0004_),
    .Q(\o_tmp[0][4] ),
    .QN(_0463_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0985_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net58),
    .D(_0011_),
    .Q(\o_tmp[0][5] ),
    .QN(_0464_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0986_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net58),
    .D(_0012_),
    .Q(\o_tmp[0][6] ),
    .QN(_0465_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0987_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net62),
    .D(_0013_),
    .Q(\o_tmp[0][7] ),
    .QN(_0466_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0988_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net62),
    .D(_0014_),
    .Q(\o_tmp[0][8] ),
    .QN(_0467_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0989_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net64),
    .D(_0015_),
    .Q(\o_tmp[0][9] ),
    .QN(_0468_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0990_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net65),
    .D(_0005_),
    .Q(\o_tmp[0][10] ),
    .QN(_0469_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0991_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net67),
    .D(_0006_),
    .Q(\o_tmp[0][11] ),
    .QN(_0470_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0992_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net69),
    .D(_0007_),
    .Q(\o_tmp[0][12] ),
    .QN(_0471_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0993_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net69),
    .D(_0008_),
    .Q(\o_tmp[0][13] ),
    .QN(_0472_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0994_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net69),
    .D(_0009_),
    .Q(\o_tmp[0][14] ),
    .QN(_0473_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0995_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net69),
    .D(_0010_),
    .Q(\o_tmp[0][15] ),
    .QN(_0474_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0996_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net50),
    .D(\o_tmp[0][0] ),
    .Q(\o_tmp[1][0] ),
    .QN(_0475_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0997_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net52),
    .D(\o_tmp[0][1] ),
    .Q(\o_tmp[1][1] ),
    .QN(_0476_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0998_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net52),
    .D(\o_tmp[0][2] ),
    .Q(\o_tmp[1][2] ),
    .QN(_0477_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _0999_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net56),
    .D(\o_tmp[0][3] ),
    .Q(\o_tmp[1][3] ),
    .QN(_0478_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1000_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net57),
    .D(\o_tmp[0][4] ),
    .Q(\o_tmp[1][4] ),
    .QN(_0479_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1001_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net58),
    .D(\o_tmp[0][5] ),
    .Q(\o_tmp[1][5] ),
    .QN(_0480_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1002_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net59),
    .D(\o_tmp[0][6] ),
    .Q(\o_tmp[1][6] ),
    .QN(_0481_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1003_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net62),
    .D(\o_tmp[0][7] ),
    .Q(\o_tmp[1][7] ),
    .QN(_0482_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1004_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net63),
    .D(\o_tmp[0][8] ),
    .Q(\o_tmp[1][8] ),
    .QN(_0483_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1005_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net64),
    .D(\o_tmp[0][9] ),
    .Q(\o_tmp[1][9] ),
    .QN(_0484_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1006_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net67),
    .D(\o_tmp[0][10] ),
    .Q(\o_tmp[1][10] ),
    .QN(_0485_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1007_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net68),
    .D(\o_tmp[0][11] ),
    .Q(\o_tmp[1][11] ),
    .QN(_0486_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1008_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net70),
    .D(\o_tmp[0][12] ),
    .Q(\o_tmp[1][12] ),
    .QN(_0487_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1009_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net70),
    .D(\o_tmp[0][13] ),
    .Q(\o_tmp[1][13] ),
    .QN(_0488_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1010_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net73),
    .D(\o_tmp[0][14] ),
    .Q(\o_tmp[1][14] ),
    .QN(_0489_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1011_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net73),
    .D(\o_tmp[0][15] ),
    .Q(\o_tmp[1][15] ),
    .QN(_0490_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1012_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net50),
    .D(\o_tmp[1][0] ),
    .Q(\o_tmp[2][0] ),
    .QN(_0491_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1013_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net53),
    .D(\o_tmp[1][1] ),
    .Q(\o_tmp[2][1] ),
    .QN(_0492_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1014_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net52),
    .D(\o_tmp[1][2] ),
    .Q(\o_tmp[2][2] ),
    .QN(_0493_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1015_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net56),
    .D(\o_tmp[1][3] ),
    .Q(\o_tmp[2][3] ),
    .QN(_0494_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1016_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net57),
    .D(\o_tmp[1][4] ),
    .Q(\o_tmp[2][4] ),
    .QN(_0495_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1017_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net58),
    .D(\o_tmp[1][5] ),
    .Q(\o_tmp[2][5] ),
    .QN(_0496_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1018_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net59),
    .D(\o_tmp[1][6] ),
    .Q(\o_tmp[2][6] ),
    .QN(_0497_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1019_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net62),
    .D(\o_tmp[1][7] ),
    .Q(\o_tmp[2][7] ),
    .QN(_0498_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1020_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net64),
    .D(\o_tmp[1][8] ),
    .Q(\o_tmp[2][8] ),
    .QN(_0499_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1021_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net65),
    .D(\o_tmp[1][9] ),
    .Q(\o_tmp[2][9] ),
    .QN(_0500_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1022_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net67),
    .D(\o_tmp[1][10] ),
    .Q(\o_tmp[2][10] ),
    .QN(_0501_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1023_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net68),
    .D(\o_tmp[1][11] ),
    .Q(\o_tmp[2][11] ),
    .QN(_0502_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1024_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net71),
    .D(\o_tmp[1][12] ),
    .Q(\o_tmp[2][12] ),
    .QN(_0503_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1025_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net71),
    .D(\o_tmp[1][13] ),
    .Q(\o_tmp[2][13] ),
    .QN(_0504_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1026_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net71),
    .D(\o_tmp[1][14] ),
    .Q(\o_tmp[2][14] ),
    .QN(_0505_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1027_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net73),
    .D(\o_tmp[1][15] ),
    .Q(\o_tmp[2][15] ),
    .QN(_0506_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1028_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net50),
    .D(\o_tmp[2][0] ),
    .Q(net34),
    .QN(_0507_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1029_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net51),
    .D(\o_tmp[2][1] ),
    .Q(net41),
    .QN(_0508_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1030_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net53),
    .D(\o_tmp[2][2] ),
    .Q(net42),
    .QN(_0509_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1031_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net56),
    .D(\o_tmp[2][3] ),
    .Q(net43),
    .QN(_0510_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1032_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net57),
    .D(\o_tmp[2][4] ),
    .Q(net44),
    .QN(_0511_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1033_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net59),
    .D(\o_tmp[2][5] ),
    .Q(net45),
    .QN(_0512_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1034_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net60),
    .D(\o_tmp[2][6] ),
    .Q(net46),
    .QN(_0513_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1035_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net63),
    .D(\o_tmp[2][7] ),
    .Q(net47),
    .QN(_0514_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1036_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net64),
    .D(\o_tmp[2][8] ),
    .Q(net48),
    .QN(_0515_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1037_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net65),
    .D(\o_tmp[2][9] ),
    .Q(net49),
    .QN(_0516_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1038_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net67),
    .D(\o_tmp[2][10] ),
    .Q(net35),
    .QN(_0517_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1039_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net68),
    .D(\o_tmp[2][11] ),
    .Q(net36),
    .QN(_0518_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1040_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net71),
    .D(\o_tmp[2][12] ),
    .Q(net37),
    .QN(_0519_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1041_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net72),
    .D(\o_tmp[2][13] ),
    .Q(net38),
    .QN(_0520_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1042_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net72),
    .D(\o_tmp[2][14] ),
    .Q(net39),
    .QN(_0521_));
 gf180mcu_osu_sc_gp9t3v3__dff_1 _1043_ (.VDD(vdd),
    .VSS(vss),
    .CLK(net73),
    .D(\o_tmp[2][15] ),
    .Q(net40),
    .QN(_0458_));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input1 (.VDD(vdd),
    .VSS(vss),
    .A(a[0]),
    .Y(net1));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input2 (.VDD(vdd),
    .VSS(vss),
    .A(a[1]),
    .Y(net2));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input3 (.VDD(vdd),
    .VSS(vss),
    .A(a[2]),
    .Y(net3));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input4 (.VDD(vdd),
    .VSS(vss),
    .A(a[3]),
    .Y(net4));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input5 (.VDD(vdd),
    .VSS(vss),
    .A(a[4]),
    .Y(net5));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input6 (.VDD(vdd),
    .VSS(vss),
    .A(a[5]),
    .Y(net6));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input7 (.VDD(vdd),
    .VSS(vss),
    .A(a[6]),
    .Y(net7));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input8 (.VDD(vdd),
    .VSS(vss),
    .A(a[7]),
    .Y(net8));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input9 (.VDD(vdd),
    .VSS(vss),
    .A(b[0]),
    .Y(net9));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input10 (.VDD(vdd),
    .VSS(vss),
    .A(b[1]),
    .Y(net10));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input11 (.VDD(vdd),
    .VSS(vss),
    .A(b[2]),
    .Y(net11));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input12 (.VDD(vdd),
    .VSS(vss),
    .A(b[3]),
    .Y(net12));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input13 (.VDD(vdd),
    .VSS(vss),
    .A(b[4]),
    .Y(net13));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input14 (.VDD(vdd),
    .VSS(vss),
    .A(b[5]),
    .Y(net14));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input15 (.VDD(vdd),
    .VSS(vss),
    .A(b[6]),
    .Y(net15));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input16 (.VDD(vdd),
    .VSS(vss),
    .A(b[7]),
    .Y(net16));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input17 (.VDD(vdd),
    .VSS(vss),
    .A(ci[0]),
    .Y(net17));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input18 (.VDD(vdd),
    .VSS(vss),
    .A(ci[10]),
    .Y(net18));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input19 (.VDD(vdd),
    .VSS(vss),
    .A(ci[11]),
    .Y(net19));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input20 (.VDD(vdd),
    .VSS(vss),
    .A(ci[12]),
    .Y(net20));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input21 (.VDD(vdd),
    .VSS(vss),
    .A(ci[13]),
    .Y(net21));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input22 (.VDD(vdd),
    .VSS(vss),
    .A(ci[14]),
    .Y(net22));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input23 (.VDD(vdd),
    .VSS(vss),
    .A(ci[15]),
    .Y(net23));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input24 (.VDD(vdd),
    .VSS(vss),
    .A(ci[1]),
    .Y(net24));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input25 (.VDD(vdd),
    .VSS(vss),
    .A(ci[2]),
    .Y(net25));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input26 (.VDD(vdd),
    .VSS(vss),
    .A(ci[3]),
    .Y(net26));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input27 (.VDD(vdd),
    .VSS(vss),
    .A(ci[4]),
    .Y(net27));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input28 (.VDD(vdd),
    .VSS(vss),
    .A(ci[5]),
    .Y(net28));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input29 (.VDD(vdd),
    .VSS(vss),
    .A(ci[6]),
    .Y(net29));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input30 (.VDD(vdd),
    .VSS(vss),
    .A(ci[7]),
    .Y(net30));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input31 (.VDD(vdd),
    .VSS(vss),
    .A(ci[8]),
    .Y(net31));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input32 (.VDD(vdd),
    .VSS(vss),
    .A(ci[9]),
    .Y(net32));
 gf180mcu_osu_sc_gp9t3v3__lshifdown input33 (.VDD(vdd),
    .VSS(vss),
    .A(clk),
    .Y(net33));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output34 (.VDD(vdd),
    .VSS(vss),
    .A(net34),
    .Y(o[0]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output35 (.VDD(vdd),
    .VSS(vss),
    .A(net35),
    .Y(o[10]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output36 (.VDD(vdd),
    .VSS(vss),
    .A(net36),
    .Y(o[11]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output37 (.VDD(vdd),
    .VSS(vss),
    .A(net37),
    .Y(o[12]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output38 (.VDD(vdd),
    .VSS(vss),
    .A(net38),
    .Y(o[13]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output39 (.VDD(vdd),
    .VSS(vss),
    .A(net39),
    .Y(o[14]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output40 (.VDD(vdd),
    .VSS(vss),
    .A(net40),
    .Y(o[15]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output41 (.VDD(vdd),
    .VSS(vss),
    .A(net41),
    .Y(o[1]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output42 (.VDD(vdd),
    .VSS(vss),
    .A(net42),
    .Y(o[2]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output43 (.VDD(vdd),
    .VSS(vss),
    .A(net43),
    .Y(o[3]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output44 (.VDD(vdd),
    .VSS(vss),
    .A(net44),
    .Y(o[4]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output45 (.VDD(vdd),
    .VSS(vss),
    .A(net45),
    .Y(o[5]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output46 (.VDD(vdd),
    .VSS(vss),
    .A(net46),
    .Y(o[6]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output47 (.VDD(vdd),
    .VSS(vss),
    .A(net47),
    .Y(o[7]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output48 (.VDD(vdd),
    .VSS(vss),
    .A(net48),
    .Y(o[8]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown output49 (.VDD(vdd),
    .VSS(vss),
    .A(net49),
    .Y(o[9]));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout50 (.VDD(vdd),
    .VSS(vss),
    .A(net55),
    .Y(net50));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout51 (.VDD(vdd),
    .VSS(vss),
    .A(net55),
    .Y(net51));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout52 (.VDD(vdd),
    .VSS(vss),
    .A(net54),
    .Y(net52));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout53 (.VDD(vdd),
    .VSS(vss),
    .A(net54),
    .Y(net53));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout54 (.VDD(vdd),
    .VSS(vss),
    .A(net55),
    .Y(net54));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout55 (.VDD(vdd),
    .VSS(vss),
    .A(net61),
    .Y(net55));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout56 (.VDD(vdd),
    .VSS(vss),
    .A(net60),
    .Y(net56));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout57 (.VDD(vdd),
    .VSS(vss),
    .A(net60),
    .Y(net57));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout58 (.VDD(vdd),
    .VSS(vss),
    .A(net59),
    .Y(net58));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout59 (.VDD(vdd),
    .VSS(vss),
    .A(net60),
    .Y(net59));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout60 (.VDD(vdd),
    .VSS(vss),
    .A(net61),
    .Y(net60));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout61 (.VDD(vdd),
    .VSS(vss),
    .A(net78),
    .Y(net61));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout62 (.VDD(vdd),
    .VSS(vss),
    .A(net66),
    .Y(net62));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout63 (.VDD(vdd),
    .VSS(vss),
    .A(net66),
    .Y(net63));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout64 (.VDD(vdd),
    .VSS(vss),
    .A(net66),
    .Y(net64));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout65 (.VDD(vdd),
    .VSS(vss),
    .A(net66),
    .Y(net65));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout66 (.VDD(vdd),
    .VSS(vss),
    .A(net77),
    .Y(net66));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout67 (.VDD(vdd),
    .VSS(vss),
    .A(net76),
    .Y(net67));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout68 (.VDD(vdd),
    .VSS(vss),
    .A(net76),
    .Y(net68));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout69 (.VDD(vdd),
    .VSS(vss),
    .A(net75),
    .Y(net69));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout70 (.VDD(vdd),
    .VSS(vss),
    .A(net75),
    .Y(net70));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout71 (.VDD(vdd),
    .VSS(vss),
    .A(net74),
    .Y(net71));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout72 (.VDD(vdd),
    .VSS(vss),
    .A(net74),
    .Y(net72));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout73 (.VDD(vdd),
    .VSS(vss),
    .A(net75),
    .Y(net73));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout74 (.VDD(vdd),
    .VSS(vss),
    .A(net75),
    .Y(net74));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout75 (.VDD(vdd),
    .VSS(vss),
    .A(net76),
    .Y(net75));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout76 (.VDD(vdd),
    .VSS(vss),
    .A(net77),
    .Y(net76));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout77 (.VDD(vdd),
    .VSS(vss),
    .A(net78),
    .Y(net77));
 gf180mcu_osu_sc_gp9t3v3__lshifdown fanout78 (.VDD(vdd),
    .VSS(vss),
    .A(net33),
    .Y(net78));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_1730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_1738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_0_1742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_2229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_2241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_2727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_2735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_2739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_3225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_3233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_0_3237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_3724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_3732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_3736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_4222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_4230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_0_4234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_4721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_4729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_4733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_5225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_0_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_5231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_5717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_0_5729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_6216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_6228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_6714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_6722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_0_6726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_7221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_7225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_7711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_7719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_7723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_8209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_8217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_0_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_8708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_0_8716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_0_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_0_8966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_0_8974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_2_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_2_8909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_2_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_2_8921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_14_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_14_8909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_14_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_14_8921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_27_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_27_8909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_27_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_27_8921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_38_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_38_4717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_38_4725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_38_4727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_38_8967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_38_8975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_39_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_39_3453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_39_3805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_39_3813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_39_3817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_39_3819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_39_3880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_39_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_39_3892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_39_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_39_4197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_39_4472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_39_4474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_39_4497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_39_4505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_39_4507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_39_4731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_39_4735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_39_5385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_39_5393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_39_8922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_40_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_40_3498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_40_3500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_40_3820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_40_3919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_40_3923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_40_4062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_40_4111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_40_4119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_40_4123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_40_4156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_40_4164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_40_4166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_40_4449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_40_4457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_40_4522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_40_4530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_40_4534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_40_4631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_40_4639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_40_4643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_40_4824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_40_5099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_40_5103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_40_5142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_40_5379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_40_5383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_40_8968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_3236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_3414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_3422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_3492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_3494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_3540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_3542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_3689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_3802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_3804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_3833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_4037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_4039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_4257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_4409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_4417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_4499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_4600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_4707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_4715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_4791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_4799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_4803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_5028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_5162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_5166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_41_5564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_5572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_5704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_41_5706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_41_8970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_41_8974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_3027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_3035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_3164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_3170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_3404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_3491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_3493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_3637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_3641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_3738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_3835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_3868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_4049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_4057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_4063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_4086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_4094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_4098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_4195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_4260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_4268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_4270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_4463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_4471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_4542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_4641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_4649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_4735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_4743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_4747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_4868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_4948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_4956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_5052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_5186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_5194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_5198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_5327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_5331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_5396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_5404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_5406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_5634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_5638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_5683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_5687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_5752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_42_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_42_5762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_5906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_6022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_42_8964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_42_8972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_2712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_2716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_2881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_3026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_3034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_3038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_3081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_3147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_3155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_3159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_3161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_3365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_3480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_3562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_3780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_3788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_3794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_3890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_3894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_4118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_4261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_4265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_4267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_4331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_4414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_4422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_4426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_4428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_4457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_4465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_4467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_4499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_4507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_4748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_4756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_4872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_4884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_4917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_5081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_5089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_5093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_5126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_5130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_5132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_5161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_5380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_5382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_5566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_5621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_5623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_5656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_5707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_5882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_6030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_6038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_6040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_6105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_6186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_43_6190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_6526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_43_8962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_43_8970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_43_8974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_2792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_2794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_3010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_3018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_3236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_3244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_3324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_3332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_3478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_3486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_3836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_3877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_3885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_3889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_3971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_3979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_3983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_4081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_4085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_4087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_4280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_4455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_4463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_4467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_4469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_4626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_4760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_4823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_4827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_4829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_4861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_4865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_4985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_4989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_4991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_5071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_5079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_5112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_5122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_5161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_5165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_5167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_5295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_5303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_5307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_5341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_5349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_5353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_5418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_5668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_5672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_5704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_5898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_6222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_6226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_6228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_44_6292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_6300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_44_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_44_6491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_44_8972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_2666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_2790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_2798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_2802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_3019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_3087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_3186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_3218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_3222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_3334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_3530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_3534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_3752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_3826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_3830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_3832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_3937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_3941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_4086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_4090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_4289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_4291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_4420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_4470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_4502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_4807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_4815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_4819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_4984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_5063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_5071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_5119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_5127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_5208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_5334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_5342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_5346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_5380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_5384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_5449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_5457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_5521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_5529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_5601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_5605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_5634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_5642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_5644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_5882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_5890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_5894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_5896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_6140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_6228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_6236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_45_6308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_6316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_45_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_45_6376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_6380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_45_8975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_1246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_1250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_1347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_1379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_1387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_1391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_2747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_2755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_2759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_2972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_2980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_2984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_2986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_3082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_3086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_3377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_3381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_3454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_3566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_3743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_3747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_3811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_3815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_4073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_4081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_4085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_4117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_4149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_4200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_4245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_4257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_4342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_4494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_4555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_4559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_4783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_5014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_5018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_5227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_5235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_5324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_5588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_5697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_5701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_5782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_5790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_5912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_5916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_6037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_6041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_6083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_6091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_6156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_46_6225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_46_6233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_46_8973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_46_8975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_1207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_1403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_2728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_2732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_3123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_3205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_3410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_3418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_3422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_3521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_3525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_3558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_3566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_4069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_4265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_4348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_4350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_4395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_4403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_4497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_4562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_4814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_5116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_5300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_5512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_5514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_5639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_5787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_5795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_5799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_5801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_5901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_5909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_5913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_6038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_47_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_6197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_6201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_6386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_47_6390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_47_6392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_47_8972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_1390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_1394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_1476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_2791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_2799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_2803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_2897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_2905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_2911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_3292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_3300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_3388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_3394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_3459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_3555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_3563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_3779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_3787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_3791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_3859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_3861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_4070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_4078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_4082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_4181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_4193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_4195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_4266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_4454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_4462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_4466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_4571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_4579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_4581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_4806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_4814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_4818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_4883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_4887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_4961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_4969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_4973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_4975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_5319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_5327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_5500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_5508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_5512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_5649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_5717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_6014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_6022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_48_6207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_6419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_48_6466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_48_8966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_48_8974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_1057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_1061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_1063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_1336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_2073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_2081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_2085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_2087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_2735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_2899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_2903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_2968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_3068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_3176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_3224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_3304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_3308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_3516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_3669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_3671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_3822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_3826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_4047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_4129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_4235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_4243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_4247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_4249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_4581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_4585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_4587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_4948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_4956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_4958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_5257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_5265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_5269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_5407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_5473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_5477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_5626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_5634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_5638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_5640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_6069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_6077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_49_6079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_6179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_6187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_6191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_49_6407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_49_6783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_6791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_49_8974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_1255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_1263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_1267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_2037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_2850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_2854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_2856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_2921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_3051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_3055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_3190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_3192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_3410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_3656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_3834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_3842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_3846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_3879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_3887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_3891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_4243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_4245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_4505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_4566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_4631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_4635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_4965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_4969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_5272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_5512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_6088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_6174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_6182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_50_6225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_6233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_6463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_50_6467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_6869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_50_8970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_50_8974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_1061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_1071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_1313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_1321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_1327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_2001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_2005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_2536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_2548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_2550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_2904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_3157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_3631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_4255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_4645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_4824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_4828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_4830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_4933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_4941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_6161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_6169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_6175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_6319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_51_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_6504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_6506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_7004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_7010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_51_8916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_51_8920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_51_8922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_52_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_52_1126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_52_1371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_1379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_1381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_2071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_2842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_3164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_52_3647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_3655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_52_3761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_3765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_4284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_4286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_52_4495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_4503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_4505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_4758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_4760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_52_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_52_4936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_4940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_4942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_52_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_5012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_52_6185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_52_6222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_6230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_52_6376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_52_6674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_6837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_52_8967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_52_8975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_1135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_1139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_1194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_1198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_1348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_1350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_2136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_2140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_2607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_2611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_2891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_2899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_3174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_3274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_3282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_3636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_3644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_3646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_4300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_4526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_4530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_4532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_4600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_4652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_4962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_4970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_5009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_5017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_5083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_5091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_5095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_53_5528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_6268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_6276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_6278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_6568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_6993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_6995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_53_8965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_53_8973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_53_8975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_1145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_2198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_2202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_2204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_2942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_2950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_2954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_2956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_3390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_3398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_3739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_3743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_3797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_4296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_4298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_4411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_4596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_4811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_4819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_5142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_5150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_5154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_5317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_5329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_5587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_5595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_5842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_6344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_6449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_6457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_6683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_6691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_6695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_6697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_6751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_54_6759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_6763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_54_7054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_7062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_54_7064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_54_8974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_55_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_2728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_55_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_3013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_55_3514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_55_3740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_3748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_55_3752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_55_3754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_55_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_3928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_55_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_4522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_55_4526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_4977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_55_4981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_55_5384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_55_5396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_55_5398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_55_5500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_55_5759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_5767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_55_5771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_55_5773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_55_6351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_55_6359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_55_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_6949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_55_6953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_55_8972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_56_4625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_56_4633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_56_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_56_4639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_56_4993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_56_5048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_56_5137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_56_5145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_56_5403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_56_5672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_56_5676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_56_5678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_56_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_56_5944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_56_5948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_56_6126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_56_6134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_56_6138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_56_6140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_56_6702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_56_6706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_56_6708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_56_6794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_56_6802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_56_6806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_56_8968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_57_8972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_63_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_63_8909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_63_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_63_8921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_75_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_75_8909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_75_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_75_8921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_87_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_87_8909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_4 FILLER_87_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_87_8921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_1397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_1407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_1957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_1967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_2517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_2527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_3077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_3085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_3087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_3637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_3645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_3647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_4197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_4205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_4207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_4757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_4765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_4767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_5317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_5325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_5327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_5877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_5885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_5887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_6437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_6445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_6447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_6997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_7005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_7007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_7557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_7565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_7567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_8117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_8125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_8127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_8677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_8685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_8687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_8965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_8973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_osu_sc_gp9t3v3__fill_1 FILLER_88_8975 (.VDD(vdd),
    .VSS(vss));
endmodule
