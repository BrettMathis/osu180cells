magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect 631 23868 5755 29130
rect 322 17407 629 19962
rect 1449 9381 1508 9422
rect 2249 9381 2303 9405
rect 3188 2700 3233 2702
<< mvpmos >>
rect 5069 27951 5189 28633
rect 5294 27951 5414 28633
rect 5069 27176 5189 27858
rect 5294 27176 5414 27858
<< mvndiff >>
rect 5543 536 5627 555
rect 5543 208 5562 536
rect 5608 208 5627 536
rect 5543 189 5627 208
<< mvpdiff >>
rect 4963 27951 5069 28633
rect 5189 27951 5294 28633
rect 5414 27951 5520 28633
rect 4963 27176 5069 27858
rect 5189 27176 5294 27858
rect 5414 27176 5520 27858
<< mvndiffc >>
rect 5562 208 5608 536
<< metal1 >>
rect 487 27093 563 27105
rect 487 27041 499 27093
rect 551 27041 563 27093
rect 487 27029 563 27041
rect 702 18378 778 18390
rect 702 18326 714 18378
rect 766 18326 778 18378
rect 702 18314 778 18326
rect 1717 18386 2025 18406
rect 1717 18334 1747 18386
rect 1799 18334 1933 18386
rect 1985 18334 2025 18386
rect 1717 18314 2025 18334
rect 2955 18386 3263 18406
rect 2955 18334 2985 18386
rect 3037 18334 3171 18386
rect 3223 18334 3263 18386
rect 2955 18314 3263 18334
rect 4194 18386 4502 18406
rect 4194 18334 4224 18386
rect 4276 18334 4410 18386
rect 4462 18334 4502 18386
rect 4194 18314 4502 18334
rect 5441 18378 5517 18390
rect 5441 18326 5453 18378
rect 5505 18326 5517 18378
rect 5441 18314 5517 18326
rect 4824 16415 5132 16435
rect 4824 16363 4854 16415
rect 4906 16363 5040 16415
rect 5092 16363 5132 16415
rect 4824 16343 5132 16363
rect 3675 16190 4437 16230
rect 3675 16138 3713 16190
rect 3765 16138 3924 16190
rect 3976 16138 4136 16190
rect 4188 16138 4347 16190
rect 4399 16138 4437 16190
rect 3675 16097 4437 16138
rect 487 15953 563 15965
rect 487 15901 499 15953
rect 551 15901 563 15953
rect 487 15889 563 15901
rect 2258 15936 2350 15977
rect 2258 15884 2278 15936
rect 2330 15884 2350 15936
rect 2258 15750 2350 15884
rect 2258 15698 2278 15750
rect 2330 15698 2350 15750
rect 2258 15658 2350 15698
rect 5344 10246 5438 11053
rect 5344 10194 5365 10246
rect 5417 10194 5438 10246
rect 5344 10076 5438 10194
rect 5345 10060 5437 10076
rect 5345 10008 5365 10060
rect 5417 10008 5437 10060
rect 5345 9967 5437 10008
rect 617 8870 925 8890
rect 617 8818 647 8870
rect 699 8818 833 8870
rect 885 8818 925 8870
rect 617 8798 925 8818
rect 2706 8739 2790 9047
rect 461 8530 553 8570
rect 461 8478 481 8530
rect 533 8478 553 8530
rect 461 8344 553 8478
rect 461 8292 481 8344
rect 533 8292 553 8344
rect 461 8251 553 8292
rect 3416 7668 3620 7806
rect 1511 6327 1603 6368
rect 1511 6275 1531 6327
rect 1583 6275 1603 6327
rect 1511 6141 1603 6275
rect 1511 6089 1531 6141
rect 1583 6089 1603 6141
rect 1511 6049 1603 6089
rect 4639 5597 4715 5609
rect 4639 5441 4651 5597
rect 4703 5441 4715 5597
rect 4639 5429 4715 5441
rect 5125 5597 5201 5609
rect 5125 5441 5137 5597
rect 5189 5441 5201 5597
rect 5125 5429 5201 5441
rect 2257 3610 2349 3650
rect 2257 3558 2277 3610
rect 2329 3558 2349 3610
rect 2257 3424 2349 3558
rect 2257 3372 2277 3424
rect 2329 3372 2349 3424
rect 2257 3331 2349 3372
rect 2397 913 2470 1034
rect 2621 913 2741 1033
rect 3346 913 3466 1033
rect 2621 376 2741 566
rect 3346 376 3466 566
rect 5547 556 5623 568
rect 5547 192 5559 556
rect 5611 192 5623 556
rect 5547 180 5623 192
rect 828 -94 1008 -82
rect 828 -146 840 -94
rect 996 -146 1008 -94
rect 828 -158 1008 -146
rect 3000 -2259 3076 -2247
rect 3000 -2415 3012 -2259
rect 3064 -2415 3076 -2259
rect 3000 -2427 3076 -2415
<< via1 >>
rect 499 27041 551 27093
rect 714 18326 766 18378
rect 1747 18334 1799 18386
rect 1933 18334 1985 18386
rect 2985 18334 3037 18386
rect 3171 18334 3223 18386
rect 4224 18334 4276 18386
rect 4410 18334 4462 18386
rect 5453 18326 5505 18378
rect 4854 16363 4906 16415
rect 5040 16363 5092 16415
rect 3713 16138 3765 16190
rect 3924 16138 3976 16190
rect 4136 16138 4188 16190
rect 4347 16138 4399 16190
rect 499 15901 551 15953
rect 2278 15884 2330 15936
rect 2278 15698 2330 15750
rect 5365 10194 5417 10246
rect 5365 10008 5417 10060
rect 647 8818 699 8870
rect 833 8818 885 8870
rect 481 8478 533 8530
rect 481 8292 533 8344
rect 1531 6275 1583 6327
rect 1531 6089 1583 6141
rect 4651 5441 4703 5597
rect 5137 5441 5189 5597
rect 2277 3558 2329 3610
rect 2277 3372 2329 3424
rect 5559 536 5611 556
rect 5559 208 5562 536
rect 5562 208 5608 536
rect 5608 208 5611 536
rect 5559 192 5611 208
rect 840 -146 996 -94
rect 3012 -2415 3064 -2259
<< metal2 >>
rect 487 27093 563 27105
rect 487 27041 499 27093
rect 551 27041 563 27093
rect 487 27029 563 27041
rect 497 15965 553 27029
rect 678 21186 772 21224
rect 678 21130 697 21186
rect 753 21130 772 21186
rect 678 21091 772 21130
rect 1732 20867 1826 20905
rect 1732 20811 1751 20867
rect 1807 20811 1826 20867
rect 1732 20772 1826 20811
rect 1916 20538 2010 20576
rect 1916 20482 1935 20538
rect 1991 20482 2010 20538
rect 1916 20443 2010 20482
rect 2970 20216 3064 20254
rect 2970 20160 2989 20216
rect 3045 20160 3064 20216
rect 2970 20121 3064 20160
rect 3155 19565 3249 19603
rect 3155 19509 3174 19565
rect 3230 19509 3249 19565
rect 3155 19470 3249 19509
rect 4209 19252 4303 19290
rect 4209 19196 4228 19252
rect 4284 19196 4303 19252
rect 4209 19157 4303 19196
rect 4393 18926 4487 18964
rect 4393 18870 4412 18926
rect 4468 18870 4487 18926
rect 4393 18831 4487 18870
rect 5447 18611 5541 18649
rect 5447 18555 5466 18611
rect 5522 18555 5541 18611
rect 5447 18516 5541 18555
rect 702 18378 778 18390
rect 702 18326 714 18378
rect 766 18326 778 18378
rect 702 16551 778 18326
rect 1717 18386 2025 18406
rect 1717 18334 1747 18386
rect 1799 18334 1933 18386
rect 1985 18334 2025 18386
rect 1717 18314 2025 18334
rect 2955 18386 3263 18406
rect 2955 18334 2985 18386
rect 3037 18334 3171 18386
rect 3223 18334 3263 18386
rect 2955 18314 3263 18334
rect 4194 18386 4502 18406
rect 4194 18334 4224 18386
rect 4276 18334 4410 18386
rect 4462 18334 4502 18386
rect 4194 18314 4502 18334
rect 5441 18378 5517 18390
rect 5441 18326 5453 18378
rect 5505 18326 5517 18378
rect 1826 16645 1916 18314
rect 3065 16645 3154 18314
rect 4303 16646 4393 18314
rect 5441 16435 5517 18326
rect 4824 16415 5517 16435
rect 4824 16363 4854 16415
rect 4906 16363 5040 16415
rect 5092 16363 5517 16415
rect 4824 16343 5517 16363
rect 3675 16192 4437 16230
rect 3675 16136 3711 16192
rect 3767 16136 3922 16192
rect 3978 16136 4134 16192
rect 4190 16136 4345 16192
rect 4401 16136 4437 16192
rect 3675 16097 4437 16136
rect 487 15953 563 15965
rect 487 15901 499 15953
rect 551 15901 563 15953
rect 487 15889 563 15901
rect 2072 10264 2166 15979
rect 2258 15945 2350 15976
rect 2256 15936 2351 15945
rect 2256 15884 2278 15936
rect 2330 15884 2351 15936
rect 2256 15750 2351 15884
rect 2256 15698 2278 15750
rect 2330 15698 2351 15750
rect 1004 10199 1913 10255
rect 831 8890 926 8894
rect 617 8870 926 8890
rect 617 8818 647 8870
rect 699 8818 833 8870
rect 885 8818 926 8870
rect 617 8798 926 8818
rect 461 8530 553 8570
rect 461 8478 481 8530
rect 533 8478 553 8530
rect 461 8434 553 8478
rect 460 8344 554 8434
rect 460 8292 481 8344
rect 533 8292 554 8344
rect 460 8 554 8292
rect 831 7826 926 8798
rect 831 7735 1156 7826
rect 1061 5893 1156 7735
rect 1857 7696 1913 10199
rect 1857 7640 2004 7696
rect 845 5795 1156 5893
rect 1508 6367 1602 6374
rect 1508 6327 1603 6367
rect 1508 6275 1531 6327
rect 1583 6275 1603 6327
rect 1508 6141 1603 6275
rect 1508 6089 1531 6141
rect 1583 6089 1603 6141
rect 1508 6049 1603 6089
rect 1948 6083 2004 7640
rect 2256 7648 2351 15698
rect 2441 12631 2535 15979
rect 2441 12575 2460 12631
rect 2516 12575 2535 12631
rect 2441 12445 2535 12575
rect 2441 12389 2460 12445
rect 2516 12389 2535 12445
rect 2441 11855 2535 12389
rect 2441 11799 2460 11855
rect 2516 11799 2535 11855
rect 2441 11669 2535 11799
rect 2441 11613 2460 11669
rect 2516 11613 2535 11669
rect 2441 10939 2535 11613
rect 2441 10883 2460 10939
rect 2516 10883 2535 10939
rect 2441 10753 2535 10883
rect 2441 10697 2460 10753
rect 2516 10697 2535 10753
rect 2441 10264 2535 10697
rect 5345 10246 5437 10286
rect 5345 10198 5365 10246
rect 5344 10194 5365 10198
rect 5417 10198 5437 10246
rect 5417 10194 5438 10198
rect 5344 10060 5438 10194
rect 5344 10008 5365 10060
rect 5417 10008 5438 10060
rect 4233 8346 4327 8525
rect 4692 8467 4786 8646
rect 4692 8370 5050 8467
rect 4233 8249 4435 8346
rect 4956 8229 5050 8370
rect 2256 7566 2859 7648
rect 845 1465 940 5795
rect 1508 5771 1602 6049
rect 1308 5647 1602 5771
rect 1877 6027 2004 6083
rect 845 1287 958 1465
rect 878 -82 958 1287
rect 1308 -1 1402 5647
rect 1877 1860 1933 6027
rect 2298 5006 2354 5866
rect 2764 5052 2859 7566
rect 4395 5916 4715 6050
rect 5344 6002 5438 10008
rect 4639 5597 4715 5916
rect 4639 5441 4651 5597
rect 4703 5441 4715 5597
rect 4639 5429 4715 5441
rect 5125 5905 5438 6002
rect 5125 5597 5201 5905
rect 5125 5441 5137 5597
rect 5189 5441 5201 5597
rect 5125 5429 5201 5441
rect 2131 4996 2354 5006
rect 2131 4940 2141 4996
rect 2301 4940 2354 4996
rect 2480 4974 2859 5052
rect 2131 4930 2311 4940
rect 2480 4655 2575 4974
rect 2256 4533 2575 4655
rect 2256 3610 2351 4533
rect 2256 3558 2277 3610
rect 2329 3558 2351 3610
rect 2256 3424 2351 3558
rect 2256 3372 2277 3424
rect 2329 3372 2351 3424
rect 2256 3331 2351 3372
rect 1877 1804 1984 1860
rect 1928 993 1984 1804
rect 1928 917 2054 993
rect 828 -94 1008 -82
rect 828 -146 840 -94
rect 996 -146 1008 -94
rect 828 -158 1008 -146
rect 1998 -1900 2054 917
rect 5547 558 5623 568
rect 5547 190 5557 558
rect 5613 190 5623 558
rect 5547 180 5623 190
rect 1998 -1956 3066 -1900
rect 3010 -2247 3066 -1956
rect 3000 -2259 3076 -2247
rect 3000 -2415 3012 -2259
rect 3064 -2415 3076 -2259
rect 3000 -2427 3076 -2415
<< via2 >>
rect 697 21130 753 21186
rect 1751 20811 1807 20867
rect 1935 20482 1991 20538
rect 2989 20160 3045 20216
rect 3174 19509 3230 19565
rect 4228 19196 4284 19252
rect 4412 18870 4468 18926
rect 5466 18555 5522 18611
rect 3711 16190 3767 16192
rect 3711 16138 3713 16190
rect 3713 16138 3765 16190
rect 3765 16138 3767 16190
rect 3711 16136 3767 16138
rect 3922 16190 3978 16192
rect 3922 16138 3924 16190
rect 3924 16138 3976 16190
rect 3976 16138 3978 16190
rect 3922 16136 3978 16138
rect 4134 16190 4190 16192
rect 4134 16138 4136 16190
rect 4136 16138 4188 16190
rect 4188 16138 4190 16190
rect 4134 16136 4190 16138
rect 4345 16190 4401 16192
rect 4345 16138 4347 16190
rect 4347 16138 4399 16190
rect 4399 16138 4401 16190
rect 4345 16136 4401 16138
rect 2460 12575 2516 12631
rect 2460 12389 2516 12445
rect 2460 11799 2516 11855
rect 2460 11613 2516 11669
rect 2460 10883 2516 10939
rect 2460 10697 2516 10753
rect 2141 4940 2301 4996
rect 5557 556 5613 558
rect 5557 192 5559 556
rect 5559 192 5611 556
rect 5611 192 5613 556
rect 5557 190 5613 192
<< metal3 >>
rect -1 21417 324 23394
rect 678 21186 772 21224
rect 678 21130 697 21186
rect 753 21130 772 21186
rect 678 21091 772 21130
rect 1732 20867 1826 20905
rect 1732 20811 1751 20867
rect 1807 20811 1826 20867
rect 1732 20772 1826 20811
rect 1916 20538 2010 20576
rect 1916 20482 1935 20538
rect 1991 20482 2010 20538
rect 1916 20443 2010 20482
rect 2970 20216 3064 20254
rect 2970 20160 2989 20216
rect 3045 20160 3064 20216
rect 2970 20121 3064 20160
rect 3155 19565 3249 19603
rect 3155 19509 3174 19565
rect 3230 19509 3249 19565
rect 3155 19470 3249 19509
rect 4209 19252 4303 19290
rect 4209 19196 4228 19252
rect 4284 19196 4303 19252
rect 4209 19157 4303 19196
rect 4393 18926 4487 18964
rect 4393 18870 4412 18926
rect 4468 18870 4487 18926
rect 4393 18831 4487 18870
rect 5447 18611 5541 18649
rect 5447 18555 5466 18611
rect 5522 18555 5541 18611
rect 5447 18516 5541 18555
rect 377 16192 5517 16235
rect 377 16136 3711 16192
rect 3767 16136 3922 16192
rect 3978 16136 4134 16192
rect 4190 16136 4345 16192
rect 4401 16136 5517 16192
rect 377 16006 5517 16136
rect 5493 12998 5794 15720
rect 2442 12631 2535 12669
rect 2442 12575 2460 12631
rect 2516 12575 2535 12631
rect 2442 12445 2535 12575
rect 2442 12389 2460 12445
rect 2516 12389 2535 12445
rect 2442 12350 2535 12389
rect 2442 11855 2535 11893
rect 2442 11799 2460 11855
rect 2516 11799 2535 11855
rect 2442 11669 2535 11799
rect 2442 11613 2460 11669
rect 2516 11613 2535 11669
rect 2442 11574 2535 11613
rect 2442 10939 2535 10977
rect 2442 10883 2460 10939
rect 2516 10883 2535 10939
rect 2442 10753 2535 10883
rect 2442 10697 2460 10753
rect 2516 10697 2535 10753
rect 2442 10658 2535 10697
rect 318 4996 2311 5012
rect 318 4940 2141 4996
rect 2301 4940 2311 4996
rect 318 4924 2311 4940
rect 5627 3135 5794 4497
rect 5547 558 5623 568
rect 5547 190 5557 558
rect 5613 190 5623 558
rect 5547 180 5623 190
rect 5636 156 5794 611
use M1_NACTIVE4310591302024_512x8m81  M1_NACTIVE4310591302024_512x8m81_0
timestamp 1669390400
transform 1 0 5585 0 1 372
box 0 0 1 1
use M2_M1$$45012012_512x8m81  M2_M1$$45012012_512x8m81_0
timestamp 1669390400
transform 1 0 2525 0 1 16164
box -803 -67 803 66
use M2_M1$$45013036_512x8m81  M2_M1$$45013036_512x8m81_0
timestamp 1669390400
transform 1 0 4056 0 1 16164
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1669390400
transform 0 -1 5163 1 0 5519
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1669390400
transform 0 -1 4677 1 0 5519
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1669390400
transform 0 -1 918 1 0 -120
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_1
timestamp 1669390400
transform 1 0 3038 0 1 -2337
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_0
timestamp 1669390400
transform 1 0 525 0 1 27067
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_1
timestamp 1669390400
transform 1 0 740 0 1 18352
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_2
timestamp 1669390400
transform 1 0 5479 0 1 18352
box 0 0 1 1
use M2_M14310591302020_512x8m81  M2_M14310591302020_512x8m81_3
timestamp 1669390400
transform 1 0 525 0 1 15927
box 0 0 1 1
use M2_M14310591302025_512x8m81  M2_M14310591302025_512x8m81_0
timestamp 1669390400
transform 1 0 5585 0 1 374
box 0 0 1 1
use M3_M2$$43370540_512x8m81  M3_M2$$43370540_512x8m81_0
timestamp 1669390400
transform 1 0 4056 0 1 16164
box 0 0 1 1
use M3_M2$$44741676_512x8m81  M3_M2$$44741676_512x8m81_0
timestamp 1669390400
transform 1 0 2525 0 1 16164
box -803 -67 803 67
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1669390400
transform 1 0 2221 0 1 4968
box 0 0 1 1
use M3_M24310591302026_512x8m81  M3_M24310591302026_512x8m81_0
timestamp 1669390400
transform 1 0 5585 0 1 374
box 0 0 1 1
use din_512x8m81  din_512x8m81_0
timestamp 1669390400
transform 1 0 323 0 1 7812
box -223 -57 2607 8999
use m2_saout01_512x8m81  m2_saout01_512x8m81_0
timestamp 1669390400
transform 1 0 686 0 1 28987
box -89 -63 4849 2153
use mux821_512x8m81  mux821_512x8m81_0
timestamp 1669390400
transform 1 0 553 0 1 16669
box -822 81 7080 12461
use outbuf_oe_512x8m81  outbuf_oe_512x8m81_0
timestamp 1669390400
transform 1 0 632 0 1 5516
box -532 -359 5177 3324
use sa_512x8m81  sa_512x8m81_0
timestamp 1669390400
transform 1 0 632 0 1 8615
box -357 -196 5034 8146
use sacntl_2_512x8m81  sacntl_2_512x8m81_0
timestamp 1669390400
transform 1 0 632 0 1 30
box -530 -24 5176 5655
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1669390400
transform 1 0 2073 0 1 12351
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1669390400
transform 1 0 2073 0 1 11575
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1669390400
transform 1 0 2073 0 1 10659
box 0 -1 93 308
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1669390400
transform -1 0 2350 0 -1 15976
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1669390400
transform -1 0 1603 0 -1 6367
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1669390400
transform 1 0 2257 0 1 3332
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1669390400
transform 1 0 5345 0 1 9968
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1669390400
transform 1 0 461 0 1 8252
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1669390400
transform 0 -1 5132 1 0 16343
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1669390400
transform 0 -1 2025 1 0 18314
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1669390400
transform 0 -1 3263 1 0 18314
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_3
timestamp 1669390400
transform 0 -1 4502 1 0 18314
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_4
timestamp 1669390400
transform 0 -1 925 1 0 8798
box 0 0 1 1
use via2_512x8m81  via2_512x8m81_0
timestamp 1669390400
transform 1 0 5448 0 1 18517
box 0 0 1 1
use via2_512x8m81  via2_512x8m81_1
timestamp 1669390400
transform 1 0 4394 0 1 18832
box 0 0 1 1
use via2_512x8m81  via2_512x8m81_2
timestamp 1669390400
transform 1 0 4210 0 1 19158
box 0 0 1 1
use via2_512x8m81  via2_512x8m81_3
timestamp 1669390400
transform 1 0 2971 0 1 20122
box 0 0 1 1
use via2_512x8m81  via2_512x8m81_4
timestamp 1669390400
transform 1 0 3156 0 1 19471
box 0 0 1 1
use via2_512x8m81  via2_512x8m81_5
timestamp 1669390400
transform 1 0 1917 0 1 20444
box 0 0 1 1
use via2_512x8m81  via2_512x8m81_6
timestamp 1669390400
transform 1 0 1733 0 1 20773
box 0 0 1 1
use via2_512x8m81  via2_512x8m81_7
timestamp 1669390400
transform 1 0 679 0 1 21092
box 0 0 1 1
use via2_x2_512x8m81  via2_x2_512x8m81_0
timestamp 1669390400
transform 1 0 2442 0 1 12351
box 0 0 1 1
use via2_x2_512x8m81  via2_x2_512x8m81_1
timestamp 1669390400
transform 1 0 2442 0 1 11575
box 0 0 1 1
use via2_x2_512x8m81  via2_x2_512x8m81_2
timestamp 1669390400
transform 1 0 2442 0 1 10659
box 0 0 1 1
use wen_wm1_512x8m81  wen_wm1_512x8m81_0
timestamp 1669390400
transform 1 0 322 0 1 -3369
box -156 -24 4946 3287
<< labels >>
rlabel metal3 s 810 18914 810 18914 4 ypass[1]
port 1 nsew
rlabel metal3 s 810 19231 810 19231 4 ypass[2]
port 2 nsew
rlabel metal3 s 810 19548 810 19548 4 ypass[3]
port 3 nsew
rlabel metal3 s 810 20204 810 20204 4 ypass[4]
port 4 nsew
rlabel metal3 s 810 20528 810 20528 4 ypass[5]
port 5 nsew
rlabel metal3 s 810 20845 810 20845 4 ypass[6]
port 6 nsew
rlabel metal3 s 810 21162 810 21162 4 ypass[7]
port 7 nsew
rlabel metal3 s 881 1467 881 1467 4 men
port 8 nsew
rlabel metal3 s 2918 1090 2918 1090 4 vss
port 9 nsew
rlabel metal3 s 2918 2179 2918 2179 4 vss
port 9 nsew
rlabel metal3 s 810 20204 810 20204 4 ypass[4]
port 4 nsew
rlabel metal3 s 3030 3831 3030 3831 4 vdd
port 10 nsew
rlabel metal3 s 2121 406 2121 406 4 vdd
port 10 nsew
rlabel metal3 s 2796 5470 2796 5470 4 vss
port 9 nsew
rlabel metal3 s 1878 11036 1878 11036 4 vss
port 9 nsew
rlabel metal3 s 810 21162 810 21162 4 ypass[7]
port 7 nsew
rlabel metal3 s 810 20845 810 20845 4 ypass[6]
port 6 nsew
rlabel metal3 s 810 20528 810 20528 4 ypass[5]
port 5 nsew
rlabel metal3 s 810 19548 810 19548 4 ypass[3]
port 3 nsew
rlabel metal3 s 810 19231 810 19231 4 ypass[2]
port 2 nsew
rlabel metal3 s 810 18914 810 18914 4 ypass[1]
port 1 nsew
rlabel metal3 s 810 18592 810 18592 4 ypass[0]
port 11 nsew
rlabel metal3 s 933 28902 933 28902 4 vdd
port 10 nsew
rlabel metal3 s 949 22015 949 22015 4 vss
port 9 nsew
rlabel metal3 s 933 18163 933 18163 4 vdd
port 10 nsew
rlabel metal3 s 973 16898 973 16898 4 vss
port 9 nsew
rlabel metal3 s 1807 13768 1807 13768 4 vdd
port 10 nsew
rlabel metal3 s 3303 7647 3303 7647 4 vdd
port 10 nsew
rlabel metal3 s 810 18592 810 18592 4 ypass[0]
port 11 nsew
flabel metal3 s 460 -586 460 -586 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 7098 460 7098 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 3309 460 3309 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 451 460 451 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 -2915 460 -2915 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 616 -1999 616 -1999 0 FreeSans 600 0 0 0 GWEN
port 13 nsew
flabel metal3 s 460 2469 460 2469 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 23368 460 23368 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 -2245 460 -2245 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 6326 460 6326 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 12529 460 12529 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 -1323 460 -1323 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 1081 460 1081 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 17115 460 17115 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 -1766 460 -1766 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 8536 460 8536 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 13222 460 13222 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 18052 460 18052 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 644 4966 644 4966 0 FreeSans 600 0 0 0 GWE
port 15 nsew
rlabel metal2 s 4862 28732 4862 28732 4 bb[1]
port 16 nsew
rlabel metal2 s 5073 28732 5073 28732 4 bb[0]
port 17 nsew
rlabel metal2 s 3832 28737 3832 28737 4 bb[2]
port 18 nsew
rlabel metal2 s 3632 28741 3632 28741 4 bb[3]
port 19 nsew
rlabel metal2 s 2593 28734 2593 28734 4 bb[4]
port 20 nsew
rlabel metal2 s 2387 28734 2387 28734 4 bb[5]
port 21 nsew
rlabel metal2 s 1155 28741 1155 28741 4 bb[7]
port 22 nsew
rlabel metal2 s 1355 28734 1355 28734 4 bb[6]
port 23 nsew
rlabel metal2 s 5499 28732 5499 28732 4 b[0]
port 24 nsew
rlabel metal2 s 4449 28732 4449 28732 4 b[1]
port 25 nsew
rlabel metal2 s 3006 28732 3006 28732 4 b[4]
port 26 nsew
rlabel metal2 s 1972 28732 1972 28732 4 b[5]
port 27 nsew
rlabel metal2 s 1770 28732 1770 28732 4 b[6]
port 28 nsew
rlabel metal2 s 736 28732 736 28732 4 b[7]
port 29 nsew
rlabel metal2 s 4251 28732 4251 28732 4 b[2]
port 30 nsew
rlabel metal2 s 3211 28732 3211 28732 4 b[3]
port 31 nsew
rlabel metal2 s 731 28732 731 28732 4 b[7]
port 29 nsew
rlabel metal2 s 488 1730 488 1730 4 datain
port 32 nsew
rlabel metal2 s 1768 28732 1768 28732 4 b[6]
port 28 nsew
rlabel metal2 s 1976 28732 1976 28732 4 b[5]
port 27 nsew
rlabel metal2 s 3004 28732 3004 28732 4 b[4]
port 26 nsew
rlabel metal2 s 3208 28732 3208 28732 4 b[3]
port 31 nsew
rlabel metal2 s 4249 28732 4249 28732 4 b[2]
port 30 nsew
rlabel metal2 s 4451 28732 4451 28732 4 b[1]
port 25 nsew
rlabel metal2 s 5497 28732 5497 28732 4 b[0]
port 24 nsew
rlabel metal2 s 1353 28734 1353 28734 4 bb[6]
port 23 nsew
rlabel metal2 s 1151 28741 1151 28741 4 bb[7]
port 22 nsew
rlabel metal2 s 2391 28734 2391 28734 4 bb[5]
port 21 nsew
rlabel metal2 s 1351 1131 1351 1131 4 q
port 33 nsew
rlabel metal2 s 2591 28734 2591 28734 4 bb[4]
port 20 nsew
rlabel metal2 s 3628 28741 3628 28741 4 bb[3]
port 19 nsew
rlabel metal2 s 3828 28737 3828 28737 4 bb[2]
port 18 nsew
rlabel metal2 s 5071 28732 5071 28732 4 bb[0]
port 17 nsew
rlabel metal2 s 4864 28732 4864 28732 4 bb[1]
port 16 nsew
rlabel metal2 s 1351 1131 1351 1131 4 q
port 33 nsew
rlabel metal1 s 993 27082 993 27082 4 pcb
port 34 nsew
rlabel metal1 s 698 8320 698 8320 4 datain
port 32 nsew
rlabel metal1 s 993 27079 993 27079 4 pcb
port 34 nsew
rlabel metal1 s 1801 15942 1801 15942 4 pcb
port 34 nsew
flabel metal1 s 722 -3358 722 -3358 0 FreeSans 600 0 0 0 WEN
port 35 nsew
<< properties >>
string FIXED_BBOX 2864 27052 2910 29928
string GDS_END 931382
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 921646
string path 14.435 135.260 14.435 149.640 
<< end >>
