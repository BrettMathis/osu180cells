magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 3446 1094
<< pwell >>
rect -86 -86 3446 453
<< mvnmos >>
rect 124 146 244 304
rect 348 146 468 304
rect 758 215 878 331
rect 926 215 1046 331
rect 1150 215 1270 331
rect 1318 215 1438 331
rect 1618 216 1738 332
rect 1842 216 1962 332
rect 2066 216 2186 332
rect 2234 216 2354 332
rect 2502 68 2622 332
rect 2870 69 2990 333
rect 3094 69 3214 333
<< mvpmos >>
rect 124 573 224 849
rect 348 573 448 849
rect 798 582 898 782
rect 946 582 1046 782
rect 1170 582 1270 782
rect 1318 582 1418 782
rect 1558 582 1658 782
rect 1842 582 1942 782
rect 2102 582 2202 782
rect 2254 582 2354 782
rect 2522 573 2622 939
rect 2870 573 2970 939
rect 3074 573 3174 939
<< mvndiff >>
rect 1538 331 1618 332
rect 36 291 124 304
rect 36 245 49 291
rect 95 245 124 291
rect 36 146 124 245
rect 244 205 348 304
rect 244 159 273 205
rect 319 159 348 205
rect 244 146 348 159
rect 468 291 556 304
rect 468 245 497 291
rect 543 245 556 291
rect 468 146 556 245
rect 628 215 758 331
rect 878 215 926 331
rect 1046 318 1150 331
rect 1046 272 1075 318
rect 1121 272 1150 318
rect 1046 215 1150 272
rect 1270 215 1318 331
rect 1438 216 1618 331
rect 1738 319 1842 332
rect 1738 273 1767 319
rect 1813 273 1842 319
rect 1738 216 1842 273
rect 1962 319 2066 332
rect 1962 273 1991 319
rect 2037 273 2066 319
rect 1962 216 2066 273
rect 2186 216 2234 332
rect 2354 221 2502 332
rect 2354 216 2427 221
rect 1438 215 1558 216
rect 628 129 698 215
rect 626 122 698 129
rect 626 76 639 122
rect 685 76 698 122
rect 626 63 698 76
rect 1498 111 1558 215
rect 1498 98 1570 111
rect 1498 52 1511 98
rect 1557 52 1570 98
rect 2414 81 2427 216
rect 2473 81 2502 221
rect 2414 68 2502 81
rect 2622 319 2710 332
rect 2622 179 2651 319
rect 2697 179 2710 319
rect 2622 68 2710 179
rect 2782 222 2870 333
rect 2782 82 2795 222
rect 2841 82 2870 222
rect 2782 69 2870 82
rect 2990 320 3094 333
rect 2990 180 3019 320
rect 3065 180 3094 320
rect 2990 69 3094 180
rect 3214 222 3302 333
rect 3214 82 3243 222
rect 3289 82 3302 222
rect 3214 69 3302 82
rect 1498 39 1570 52
<< mvpdiff >>
rect 666 928 738 941
rect 36 836 124 849
rect 36 696 49 836
rect 95 696 124 836
rect 36 573 124 696
rect 224 836 348 849
rect 224 790 253 836
rect 299 790 348 836
rect 224 573 348 790
rect 448 632 536 849
rect 448 586 477 632
rect 523 586 536 632
rect 448 573 536 586
rect 666 788 679 928
rect 725 788 738 928
rect 2434 926 2522 939
rect 666 782 738 788
rect 2434 786 2447 926
rect 2493 786 2522 926
rect 2434 782 2522 786
rect 666 582 798 782
rect 898 582 946 782
rect 1046 735 1170 782
rect 1046 595 1075 735
rect 1121 595 1170 735
rect 1046 582 1170 595
rect 1270 582 1318 782
rect 1418 769 1558 782
rect 1418 629 1447 769
rect 1493 629 1558 769
rect 1418 582 1558 629
rect 1658 735 1842 782
rect 1658 595 1767 735
rect 1813 595 1842 735
rect 1658 582 1842 595
rect 1942 735 2102 782
rect 1942 595 1991 735
rect 2037 595 2102 735
rect 1942 582 2102 595
rect 2202 582 2254 782
rect 2354 582 2522 782
rect 2442 573 2522 582
rect 2622 726 2710 939
rect 2622 586 2651 726
rect 2697 586 2710 726
rect 2622 573 2710 586
rect 2782 926 2870 939
rect 2782 786 2795 926
rect 2841 786 2870 926
rect 2782 573 2870 786
rect 2970 726 3074 939
rect 2970 586 2999 726
rect 3045 586 3074 726
rect 2970 573 3074 586
rect 3174 926 3262 939
rect 3174 786 3203 926
rect 3249 786 3262 926
rect 3174 573 3262 786
<< mvndiffc >>
rect 49 245 95 291
rect 273 159 319 205
rect 497 245 543 291
rect 1075 272 1121 318
rect 1767 273 1813 319
rect 1991 273 2037 319
rect 639 76 685 122
rect 1511 52 1557 98
rect 2427 81 2473 221
rect 2651 179 2697 319
rect 2795 82 2841 222
rect 3019 180 3065 320
rect 3243 82 3289 222
<< mvpdiffc >>
rect 49 696 95 836
rect 253 790 299 836
rect 477 586 523 632
rect 679 788 725 928
rect 2447 786 2493 926
rect 1075 595 1121 735
rect 1447 629 1493 769
rect 1767 595 1813 735
rect 1991 595 2037 735
rect 2651 586 2697 726
rect 2795 786 2841 926
rect 2999 586 3045 726
rect 3203 786 3249 926
<< polysilicon >>
rect 2522 939 2622 983
rect 2870 939 2970 983
rect 3074 939 3174 983
rect 124 849 224 893
rect 348 849 448 893
rect 1170 874 1942 914
rect 1170 861 1270 874
rect 798 782 898 826
rect 946 782 1046 826
rect 1170 815 1183 861
rect 1229 815 1270 861
rect 1170 782 1270 815
rect 1318 782 1418 826
rect 1558 782 1658 826
rect 1842 782 1942 874
rect 2102 782 2202 826
rect 2254 782 2354 826
rect 124 400 224 573
rect 124 354 137 400
rect 183 354 224 400
rect 124 348 224 354
rect 348 431 448 573
rect 798 549 898 582
rect 798 503 811 549
rect 857 503 898 549
rect 798 490 898 503
rect 348 391 878 431
rect 348 383 468 391
rect 124 304 244 348
rect 348 337 361 383
rect 407 337 468 383
rect 348 304 468 337
rect 758 331 878 391
rect 946 410 1046 582
rect 1170 538 1270 582
rect 946 375 959 410
rect 926 364 959 375
rect 1005 364 1046 410
rect 1318 410 1418 582
rect 1558 549 1658 582
rect 1558 503 1571 549
rect 1617 503 1658 549
rect 1558 490 1658 503
rect 926 331 1046 364
rect 1150 331 1270 375
rect 1318 364 1331 410
rect 1377 375 1418 410
rect 1618 376 1658 490
rect 1842 522 1942 582
rect 2102 549 2202 582
rect 2102 538 2143 549
rect 1842 482 2038 522
rect 2130 503 2143 538
rect 2189 503 2202 549
rect 2130 490 2202 503
rect 1998 448 2038 482
rect 1998 408 2106 448
rect 2066 376 2106 408
rect 2254 411 2354 582
rect 2254 376 2295 411
rect 1377 364 1438 375
rect 1318 331 1438 364
rect 1618 332 1738 376
rect 1842 332 1962 376
rect 2066 332 2186 376
rect 2234 365 2295 376
rect 2341 365 2354 411
rect 2522 540 2622 573
rect 2522 494 2535 540
rect 2581 494 2622 540
rect 2522 376 2622 494
rect 2234 332 2354 365
rect 2502 332 2622 376
rect 2870 456 2970 573
rect 3074 456 3174 573
rect 2870 412 3174 456
rect 2870 366 2883 412
rect 2929 393 3174 412
rect 2929 366 2990 393
rect 2870 333 2990 366
rect 3094 377 3174 393
rect 3094 333 3214 377
rect 124 102 244 146
rect 348 102 468 146
rect 758 171 878 215
rect 926 171 1046 215
rect 1150 182 1270 215
rect 1150 136 1163 182
rect 1209 136 1270 182
rect 1318 171 1438 215
rect 1150 123 1270 136
rect 1618 172 1738 216
rect 1842 183 1962 216
rect 1842 137 1855 183
rect 1901 137 1962 183
rect 2066 172 2186 216
rect 2234 172 2354 216
rect 1842 124 1962 137
rect 2502 24 2622 68
rect 2870 25 2990 69
rect 3094 25 3214 69
<< polycontact >>
rect 1183 815 1229 861
rect 137 354 183 400
rect 811 503 857 549
rect 361 337 407 383
rect 959 364 1005 410
rect 1571 503 1617 549
rect 1331 364 1377 410
rect 2143 503 2189 549
rect 2295 365 2341 411
rect 2535 494 2581 540
rect 2883 366 2929 412
rect 1163 136 1209 182
rect 1855 137 1901 183
<< metal1 >>
rect 0 928 3360 1098
rect 0 918 679 928
rect 49 836 95 847
rect 242 836 310 918
rect 242 790 253 836
rect 299 790 310 836
rect 725 926 3360 928
rect 725 918 2447 926
rect 679 777 725 788
rect 771 861 1229 872
rect 771 815 1183 861
rect 771 804 1229 815
rect 95 731 660 735
rect 771 731 817 804
rect 1447 769 1493 918
rect 2493 918 2795 926
rect 2447 775 2493 786
rect 2841 918 3203 926
rect 2795 775 2841 786
rect 3249 918 3360 926
rect 3203 775 3249 786
rect 95 696 817 731
rect 49 689 817 696
rect 49 685 407 689
rect 641 685 817 689
rect 1075 735 1121 746
rect 126 400 298 430
rect 126 354 137 400
rect 183 354 298 400
rect 361 383 407 685
rect 361 308 407 337
rect 49 291 407 308
rect 95 262 407 291
rect 477 632 523 643
rect 477 560 523 586
rect 1447 618 1493 629
rect 1767 735 1813 746
rect 1075 560 1121 595
rect 477 549 857 560
rect 477 514 811 549
rect 477 291 543 514
rect 49 234 95 245
rect 477 245 497 291
rect 477 234 543 245
rect 273 205 319 216
rect 273 133 319 159
rect 811 196 857 503
rect 1075 549 1617 560
rect 1075 503 1571 549
rect 1075 492 1617 503
rect 926 364 959 410
rect 1005 364 1016 410
rect 926 242 1016 364
rect 1075 318 1121 492
rect 1767 421 1813 595
rect 1331 410 1813 421
rect 1377 364 1813 410
rect 1331 353 1813 364
rect 1075 261 1121 272
rect 1767 319 1813 353
rect 1767 262 1813 273
rect 1991 735 2411 746
rect 2037 700 2411 735
rect 1991 319 2037 595
rect 1991 262 2037 273
rect 2143 549 2189 560
rect 2143 201 2189 503
rect 2365 540 2411 700
rect 2651 726 2697 737
rect 2365 494 2535 540
rect 2581 494 2592 540
rect 2651 422 2697 586
rect 2295 412 2697 422
rect 2999 726 3065 737
rect 3045 586 3065 726
rect 2295 411 2883 412
rect 2341 366 2883 411
rect 2929 366 2940 412
rect 2341 365 2697 366
rect 2295 354 2697 365
rect 2651 319 2697 354
rect 1199 196 2189 201
rect 811 183 2189 196
rect 811 182 1855 183
rect 811 136 1163 182
rect 1209 155 1855 182
rect 1209 136 1220 155
rect 1844 137 1855 155
rect 1901 137 2189 183
rect 2427 221 2473 232
rect 273 122 685 133
rect 273 90 639 122
rect 0 76 639 90
rect 1511 98 1557 109
rect 685 76 1511 90
rect 0 52 1511 76
rect 1557 81 2427 90
rect 2999 320 3065 586
rect 2999 318 3019 320
rect 2942 242 3019 318
rect 2651 168 2697 179
rect 2795 222 2841 233
rect 2473 82 2795 90
rect 3019 169 3065 180
rect 3243 222 3289 233
rect 2841 82 3243 90
rect 3289 82 3360 90
rect 2473 81 3360 82
rect 1557 52 3360 81
rect 0 -90 3360 52
<< labels >>
flabel metal1 s 126 354 298 430 0 FreeSans 200 0 0 0 CLK
port 2 nsew clock input
flabel metal1 s 926 242 1016 410 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 2999 318 3065 737 0 FreeSans 200 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 918 3360 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 3243 232 3289 233 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2942 242 3065 318 1 Q
port 3 nsew default output
rlabel metal1 s 3019 169 3065 242 1 Q
port 3 nsew default output
rlabel metal1 s 3203 790 3249 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2795 790 2841 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2447 790 2493 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1447 790 1493 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 679 790 725 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 242 790 310 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3203 777 3249 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2795 777 2841 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2447 777 2493 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1447 777 1493 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 679 777 725 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3203 775 3249 777 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2795 775 2841 777 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2447 775 2493 777 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1447 775 1493 777 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1447 618 1493 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2795 232 2841 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3243 216 3289 232 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2795 216 2841 232 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2427 216 2473 232 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3243 133 3289 216 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2795 133 2841 216 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2427 133 2473 216 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 133 319 216 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3243 109 3289 133 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2795 109 2841 133 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2427 109 2473 133 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 109 685 133 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3243 90 3289 109 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2795 90 2841 109 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2427 90 2473 109 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1511 90 1557 109 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 90 685 109 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3360 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3360 1008
string GDS_END 584480
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 576570
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
