magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 2326 1094
<< pwell >>
rect -86 -86 2326 453
<< mvnmos >>
rect 124 92 244 250
rect 384 110 504 250
rect 752 107 872 247
rect 920 107 1040 247
rect 1144 107 1264 247
rect 1404 107 1524 265
rect 1628 107 1748 265
rect 1996 69 2116 333
<< mvpmos >>
rect 144 573 244 849
rect 404 649 504 849
rect 772 652 872 852
rect 920 652 1020 852
rect 1124 652 1224 852
rect 1364 576 1464 852
rect 1568 576 1668 852
rect 1996 573 2096 939
<< mvndiff >>
rect 36 193 124 250
rect 36 147 49 193
rect 95 147 124 193
rect 36 92 124 147
rect 244 168 384 250
rect 244 122 273 168
rect 319 122 384 168
rect 244 110 384 122
rect 504 193 592 250
rect 1908 287 1996 333
rect 1324 247 1404 265
rect 504 147 533 193
rect 579 147 592 193
rect 504 110 592 147
rect 664 193 752 247
rect 664 147 677 193
rect 723 147 752 193
rect 244 92 324 110
rect 664 107 752 147
rect 872 107 920 247
rect 1040 234 1144 247
rect 1040 188 1069 234
rect 1115 188 1144 234
rect 1040 107 1144 188
rect 1264 107 1404 247
rect 1524 166 1628 265
rect 1524 120 1553 166
rect 1599 120 1628 166
rect 1524 107 1628 120
rect 1748 252 1836 265
rect 1748 206 1777 252
rect 1823 206 1836 252
rect 1748 107 1836 206
rect 1908 147 1921 287
rect 1967 147 1996 287
rect 1908 69 1996 147
rect 2116 287 2204 333
rect 2116 147 2145 287
rect 2191 147 2204 287
rect 2116 69 2204 147
<< mvpdiff >>
rect 56 805 144 849
rect 56 665 69 805
rect 115 665 144 805
rect 56 573 144 665
rect 244 805 404 849
rect 244 665 273 805
rect 319 665 404 805
rect 244 649 404 665
rect 504 805 592 849
rect 504 665 533 805
rect 579 665 592 805
rect 504 649 592 665
rect 684 805 772 852
rect 684 665 697 805
rect 743 665 772 805
rect 684 652 772 665
rect 872 652 920 852
rect 1020 805 1124 852
rect 1020 665 1049 805
rect 1095 665 1124 805
rect 1020 652 1124 665
rect 1224 652 1364 852
rect 244 573 324 649
rect 1284 576 1364 652
rect 1464 805 1568 852
rect 1464 665 1493 805
rect 1539 665 1568 805
rect 1464 576 1568 665
rect 1668 805 1756 852
rect 1668 665 1697 805
rect 1743 665 1756 805
rect 1668 576 1756 665
rect 1908 805 1996 939
rect 1908 665 1921 805
rect 1967 665 1996 805
rect 1908 573 1996 665
rect 2096 805 2184 939
rect 2096 665 2125 805
rect 2171 665 2184 805
rect 2096 573 2184 665
<< mvndiffc >>
rect 49 147 95 193
rect 273 122 319 168
rect 533 147 579 193
rect 677 147 723 193
rect 1069 188 1115 234
rect 1553 120 1599 166
rect 1777 206 1823 252
rect 1921 147 1967 287
rect 2145 147 2191 287
<< mvpdiffc >>
rect 69 665 115 805
rect 273 665 319 805
rect 533 665 579 805
rect 697 665 743 805
rect 1049 665 1095 805
rect 1493 665 1539 805
rect 1697 665 1743 805
rect 1921 665 1967 805
rect 2125 665 2171 805
<< polysilicon >>
rect 404 944 1020 984
rect 144 849 244 893
rect 404 849 504 944
rect 772 852 872 896
rect 920 852 1020 944
rect 1996 939 2096 983
rect 1124 852 1224 896
rect 1364 852 1464 896
rect 1568 852 1668 896
rect 144 372 244 573
rect 144 326 157 372
rect 203 326 244 372
rect 144 294 244 326
rect 404 372 504 649
rect 404 326 417 372
rect 463 326 504 372
rect 404 294 504 326
rect 124 250 244 294
rect 384 250 504 294
rect 772 372 872 652
rect 920 472 1020 652
rect 1124 608 1224 652
rect 1124 592 1223 608
rect 1092 579 1223 592
rect 1092 533 1105 579
rect 1151 533 1223 579
rect 1092 520 1223 533
rect 1364 532 1464 576
rect 1568 532 1668 576
rect 920 433 1264 472
rect 1011 432 1264 433
rect 772 326 813 372
rect 859 326 872 372
rect 772 291 872 326
rect 752 247 872 291
rect 920 372 992 385
rect 920 326 933 372
rect 979 343 992 372
rect 979 326 1040 343
rect 920 247 1040 326
rect 1144 247 1264 432
rect 1404 385 1464 532
rect 1628 465 1668 532
rect 1996 465 2096 573
rect 1628 393 2096 465
rect 1404 372 1524 385
rect 1404 326 1417 372
rect 1463 326 1524 372
rect 1404 265 1524 326
rect 1628 372 1748 393
rect 1628 326 1641 372
rect 1687 326 1748 372
rect 1996 377 2096 393
rect 1996 333 2116 377
rect 1628 265 1748 326
rect 124 48 244 92
rect 384 66 504 110
rect 752 63 872 107
rect 920 63 1040 107
rect 1144 63 1264 107
rect 1404 63 1524 107
rect 1628 63 1748 107
rect 1996 25 2116 69
<< polycontact >>
rect 157 326 203 372
rect 417 326 463 372
rect 1105 533 1151 579
rect 813 326 859 372
rect 933 326 979 372
rect 1417 326 1463 372
rect 1641 326 1687 372
<< metal1 >>
rect 0 918 2240 1098
rect 49 805 115 816
rect 49 665 69 805
rect 49 654 115 665
rect 273 805 319 918
rect 273 654 319 665
rect 533 805 579 816
rect 49 269 95 654
rect 142 372 203 542
rect 533 522 579 665
rect 697 805 743 918
rect 697 654 743 665
rect 1049 805 1095 816
rect 1493 805 1539 918
rect 1095 665 1243 682
rect 1049 636 1243 665
rect 1493 654 1539 665
rect 1697 805 1747 816
rect 1743 665 1747 805
rect 1105 579 1151 590
rect 1105 522 1151 533
rect 533 476 1151 522
rect 142 326 157 372
rect 142 315 203 326
rect 417 372 463 383
rect 417 271 463 326
rect 217 269 463 271
rect 49 225 463 269
rect 49 223 231 225
rect 49 193 95 223
rect 533 193 579 476
rect 813 372 866 430
rect 859 326 866 372
rect 813 242 866 326
rect 933 372 979 476
rect 933 315 979 326
rect 1197 269 1243 636
rect 1697 475 1747 665
rect 1417 473 1747 475
rect 1921 805 1986 816
rect 1967 665 1986 805
rect 1417 429 1823 473
rect 1417 372 1463 429
rect 1417 315 1463 326
rect 1641 372 1687 383
rect 1641 269 1687 326
rect 1197 245 1687 269
rect 1069 234 1687 245
rect 49 136 95 147
rect 273 168 319 179
rect 533 136 579 147
rect 677 193 723 204
rect 1115 223 1687 234
rect 1733 252 1823 429
rect 1115 188 1238 223
rect 1733 206 1777 252
rect 1733 195 1823 206
rect 1921 287 1986 665
rect 2125 805 2171 918
rect 2125 654 2171 665
rect 1069 177 1238 188
rect 273 90 319 122
rect 677 90 723 147
rect 1553 166 1599 177
rect 1967 147 1986 287
rect 1921 136 1986 147
rect 2145 287 2191 298
rect 1553 90 1599 120
rect 2145 90 2191 147
rect 0 -90 2240 90
<< labels >>
flabel metal1 s 813 242 866 430 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 142 315 203 542 0 FreeSans 200 0 0 0 E
port 2 nsew clock input
flabel metal1 s 1921 136 1986 816 0 FreeSans 200 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 918 2240 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 2145 204 2191 298 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2125 654 2171 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1493 654 1539 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 697 654 743 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 654 319 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2145 179 2191 204 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 179 723 204 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2145 177 2191 179 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 177 723 179 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 177 319 179 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2145 90 2191 177 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 90 1599 177 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 90 723 177 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 177 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2240 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2240 1008
string GDS_END 969962
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 964198
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
