magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -80 1003 80 1062
rect -80 957 -23 1003
rect 23 957 80 1003
rect -80 839 80 957
rect -80 793 -23 839
rect 23 793 80 839
rect -80 676 80 793
rect -80 630 -23 676
rect 23 630 80 676
rect -80 513 80 630
rect -80 467 -23 513
rect 23 467 80 513
rect -80 350 80 467
rect -80 304 -23 350
rect 23 304 80 350
rect -80 186 80 304
rect -80 140 -23 186
rect 23 140 80 186
rect -80 23 80 140
rect -80 -23 -23 23
rect 23 -23 80 23
rect -80 -140 80 -23
rect -80 -186 -23 -140
rect 23 -186 80 -140
rect -80 -304 80 -186
rect -80 -350 -23 -304
rect 23 -350 80 -304
rect -80 -467 80 -350
rect -80 -513 -23 -467
rect 23 -513 80 -467
rect -80 -630 80 -513
rect -80 -676 -23 -630
rect 23 -676 80 -630
rect -80 -793 80 -676
rect -80 -839 -23 -793
rect 23 -839 80 -793
rect -80 -957 80 -839
rect -80 -1003 -23 -957
rect 23 -1003 80 -957
rect -80 -1061 80 -1003
<< psubdiffcont >>
rect -23 957 23 1003
rect -23 793 23 839
rect -23 630 23 676
rect -23 467 23 513
rect -23 304 23 350
rect -23 140 23 186
rect -23 -23 23 23
rect -23 -186 23 -140
rect -23 -350 23 -304
rect -23 -513 23 -467
rect -23 -676 23 -630
rect -23 -839 23 -793
rect -23 -1003 23 -957
<< metal1 >>
rect -71 1003 71 1053
rect -71 957 -23 1003
rect 23 957 71 1003
rect -71 839 71 957
rect -71 793 -23 839
rect 23 793 71 839
rect -71 676 71 793
rect -71 630 -23 676
rect 23 630 71 676
rect -71 513 71 630
rect -71 467 -23 513
rect 23 467 71 513
rect -71 350 71 467
rect -71 304 -23 350
rect 23 304 71 350
rect -71 186 71 304
rect -71 140 -23 186
rect 23 140 71 186
rect -71 23 71 140
rect -71 -23 -23 23
rect 23 -23 71 23
rect -71 -140 71 -23
rect -71 -186 -23 -140
rect 23 -186 71 -140
rect -71 -304 71 -186
rect -71 -350 -23 -304
rect 23 -350 71 -304
rect -71 -467 71 -350
rect -71 -513 -23 -467
rect 23 -513 71 -467
rect -71 -630 71 -513
rect -71 -676 -23 -630
rect 23 -676 71 -630
rect -71 -793 71 -676
rect -71 -839 -23 -793
rect 23 -839 71 -793
rect -71 -957 71 -839
rect -71 -1003 -23 -957
rect 23 -1003 71 -957
rect -71 -1053 71 -1003
<< properties >>
string GDS_END 226354
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 225326
<< end >>
