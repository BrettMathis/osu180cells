magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 454
rect 224 0 344 454
rect 448 0 568 454
<< mvndiff >>
rect -88 441 0 454
rect -88 395 -75 441
rect -29 395 0 441
rect -88 314 0 395
rect -88 268 -75 314
rect -29 268 0 314
rect -88 187 0 268
rect -88 141 -75 187
rect -29 141 0 187
rect -88 59 0 141
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 441 224 454
rect 120 395 149 441
rect 195 395 224 441
rect 120 314 224 395
rect 120 268 149 314
rect 195 268 224 314
rect 120 187 224 268
rect 120 141 149 187
rect 195 141 224 187
rect 120 59 224 141
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 441 448 454
rect 344 395 373 441
rect 419 395 448 441
rect 344 314 448 395
rect 344 268 373 314
rect 419 268 448 314
rect 344 187 448 268
rect 344 141 373 187
rect 419 141 448 187
rect 344 59 448 141
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 441 656 454
rect 568 395 597 441
rect 643 395 656 441
rect 568 314 656 395
rect 568 268 597 314
rect 643 268 656 314
rect 568 187 656 268
rect 568 141 597 187
rect 643 141 656 187
rect 568 59 656 141
rect 568 13 597 59
rect 643 13 656 59
rect 568 0 656 13
<< mvndiffc >>
rect -75 395 -29 441
rect -75 268 -29 314
rect -75 141 -29 187
rect -75 13 -29 59
rect 149 395 195 441
rect 149 268 195 314
rect 149 141 195 187
rect 149 13 195 59
rect 373 395 419 441
rect 373 268 419 314
rect 373 141 419 187
rect 373 13 419 59
rect 597 395 643 441
rect 597 268 643 314
rect 597 141 643 187
rect 597 13 643 59
<< polysilicon >>
rect 0 454 120 498
rect 224 454 344 498
rect 448 454 568 498
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
<< metal1 >>
rect -75 441 -29 454
rect -75 314 -29 395
rect -75 187 -29 268
rect -75 59 -29 141
rect -75 0 -29 13
rect 149 441 195 454
rect 149 314 195 395
rect 149 187 195 268
rect 149 59 195 141
rect 149 0 195 13
rect 373 441 419 454
rect 373 314 419 395
rect 373 187 419 268
rect 373 59 419 141
rect 373 0 419 13
rect 597 441 643 454
rect 597 314 643 395
rect 597 187 643 268
rect 597 59 643 141
rect 597 0 643 13
<< labels >>
flabel metal1 s -52 227 -52 227 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 227 620 227 0 FreeSans 200 0 0 0 D
flabel metal1 s 172 227 172 227 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 227 396 227 0 FreeSans 200 0 0 0 S
<< properties >>
string GDS_END 268366
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 265682
<< end >>
