magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< obsv1 >>
rect 0 0 86372 96976
<< obsv2 >>
rect 0 0 86372 96976
<< metal3 >>
rect 1401 96176 2401 96976
rect 2626 96368 3626 96976
rect 4137 96176 5137 96976
rect 5362 96368 6362 96976
rect 6801 96176 7801 96976
rect 8026 96368 9026 96976
rect 9537 96176 10537 96976
rect 10762 96368 11762 96976
rect 12201 96176 13201 96976
rect 13426 96368 14426 96976
rect 14937 96176 15937 96976
rect 16162 96368 17162 96976
rect 17601 96176 18601 96976
rect 18826 96368 19826 96976
rect 20653 96176 21653 96976
rect 22258 96368 23258 96976
rect 23483 96176 24483 96976
rect 25158 96368 26158 96976
rect 26572 96176 27572 96976
rect 27877 96368 28877 96976
rect 29273 96368 30273 96976
rect 30710 96176 31710 96976
rect 32381 96368 33381 96976
rect 34024 96368 35024 96976
rect 35415 96176 36415 96976
rect 36948 96368 37948 96976
rect 38585 96176 39585 96976
rect 39882 96368 40882 96976
rect 41230 96176 42230 96976
rect 42430 96368 43430 96976
rect 43713 96368 44713 96976
rect 45069 96176 46069 96976
rect 46313 96176 47313 96976
rect 47538 96368 48538 96976
rect 48901 96176 49901 96976
rect 50465 96368 51465 96976
rect 52569 96176 53569 96976
rect 54262 96176 55262 96976
rect 55990 96368 56990 96976
rect 57547 96176 58547 96976
rect 58791 96368 59791 96976
rect 60977 96176 61977 96976
rect 62202 96368 63202 96976
rect 63713 96176 64713 96976
rect 64938 96368 65938 96976
rect 66377 96176 67377 96976
rect 67602 96368 68602 96976
rect 69113 96176 70113 96976
rect 70338 96368 71338 96976
rect 71777 96176 72777 96976
rect 73002 96368 74002 96976
rect 74513 96176 75513 96976
rect 75738 96368 76738 96976
rect 77177 96176 78177 96976
rect 78402 96368 79402 96976
rect 80229 96176 81229 96976
rect 81834 96368 82834 96976
rect 83059 96176 84059 96976
rect 84666 96176 85666 96976
rect 0 95176 86372 96176
rect 0 94776 1014 94976
rect 25376 94776 25948 94785
rect 58855 94776 59427 94785
rect 85358 94776 86372 94976
rect 0 94728 27272 94776
rect 58855 94728 86372 94776
rect 0 94527 86372 94728
rect 0 94476 27272 94527
rect 30402 94526 54622 94527
rect 58855 94476 86372 94527
rect 0 94276 1014 94476
rect 25376 94461 25948 94476
rect 58855 94461 59427 94476
rect 85358 94276 86372 94476
rect 0 93376 1706 94076
rect 84666 93376 86372 94076
rect 0 92976 1014 93176
rect 85358 92976 86372 93176
rect 0 92928 27272 92976
rect 59421 92928 86372 92976
rect 0 92727 86372 92928
rect 0 92676 27272 92727
rect 30403 92726 54622 92727
rect 59421 92676 86372 92727
rect 0 92476 1014 92676
rect 85358 92476 86372 92676
rect 0 91576 1706 92276
rect 84666 91576 86372 92276
rect 0 91176 1014 91376
rect 85358 91176 86372 91376
rect 0 91128 27272 91176
rect 59421 91128 86372 91176
rect 0 90927 86372 91128
rect 0 90876 27272 90927
rect 30403 90926 54622 90927
rect 59421 90876 86372 90927
rect 0 90676 1014 90876
rect 85358 90676 86372 90876
rect 0 89776 1706 90476
rect 84666 89776 86372 90476
rect 0 89376 1014 89576
rect 85358 89376 86372 89576
rect 0 89328 27272 89376
rect 59421 89328 86372 89376
rect 0 89127 86372 89328
rect 0 89076 27272 89127
rect 30403 89126 54622 89127
rect 59421 89076 86372 89127
rect 0 88876 1014 89076
rect 85358 88876 86372 89076
rect 0 87976 1706 88676
rect 84666 87976 86372 88676
rect 0 87576 1014 87776
rect 85358 87576 86372 87776
rect 0 87528 27272 87576
rect 59421 87528 86372 87576
rect 0 87327 86372 87528
rect 0 87276 27272 87327
rect 30403 87326 54622 87327
rect 59421 87276 86372 87327
rect 0 87076 1014 87276
rect 85358 87076 86372 87276
rect 0 86176 1706 86876
rect 84666 86176 86372 86876
rect 0 85776 1014 85976
rect 85358 85776 86372 85976
rect 0 85728 27272 85776
rect 59421 85728 86372 85776
rect 0 85527 86372 85728
rect 0 85476 27272 85527
rect 30403 85526 54622 85527
rect 59421 85476 86372 85527
rect 0 85276 1014 85476
rect 85358 85276 86372 85476
rect 0 84376 1706 85076
rect 84666 84376 86372 85076
rect 0 83976 1014 84176
rect 85358 83976 86372 84176
rect 0 83928 27272 83976
rect 59421 83928 86372 83976
rect 0 83727 86372 83928
rect 0 83676 27272 83727
rect 30403 83726 54622 83727
rect 59421 83676 86372 83727
rect 0 83476 1014 83676
rect 85358 83476 86372 83676
rect 0 82576 1706 83276
rect 84666 82576 86372 83276
rect 0 82176 1014 82376
rect 85358 82176 86372 82376
rect 0 82128 27272 82176
rect 59421 82128 86372 82176
rect 0 81927 86372 82128
rect 0 81876 27272 81927
rect 30403 81926 54622 81927
rect 59421 81876 86372 81927
rect 0 81676 1014 81876
rect 85358 81676 86372 81876
rect 0 80776 1706 81476
rect 84666 80776 86372 81476
rect 0 80376 1014 80576
rect 85358 80376 86372 80576
rect 0 80328 27272 80376
rect 59421 80328 86372 80376
rect 0 80127 86372 80328
rect 0 80076 27272 80127
rect 30403 80126 54622 80127
rect 59421 80076 86372 80127
rect 0 79876 1014 80076
rect 85358 79876 86372 80076
rect 0 78976 1706 79676
rect 84666 78976 86372 79676
rect 0 78576 1014 78776
rect 85358 78576 86372 78776
rect 0 78528 27272 78576
rect 59421 78528 86372 78576
rect 0 78327 86372 78528
rect 0 78276 27272 78327
rect 30403 78326 54622 78327
rect 59421 78276 86372 78327
rect 0 78076 1014 78276
rect 85358 78076 86372 78276
rect 0 77176 1706 77876
rect 84666 77176 86372 77876
rect 0 76776 1014 76976
rect 85358 76776 86372 76976
rect 0 76728 27272 76776
rect 59421 76728 86372 76776
rect 0 76527 86372 76728
rect 0 76476 27272 76527
rect 30403 76526 54622 76527
rect 59421 76476 86372 76527
rect 0 76276 1014 76476
rect 85358 76276 86372 76476
rect 0 75376 1706 76076
rect 84666 75376 86372 76076
rect 0 74976 1014 75176
rect 85358 74976 86372 75176
rect 0 74928 27272 74976
rect 59421 74928 86372 74976
rect 0 74727 86372 74928
rect 0 74676 27272 74727
rect 30403 74726 54622 74727
rect 59421 74676 86372 74727
rect 0 74476 1014 74676
rect 85358 74476 86372 74676
rect 0 73576 1706 74276
rect 84666 73576 86372 74276
rect 0 73176 1014 73376
rect 85358 73176 86372 73376
rect 0 73128 27272 73176
rect 59421 73128 86372 73176
rect 0 72927 86372 73128
rect 0 72876 27272 72927
rect 30403 72926 54622 72927
rect 59421 72876 86372 72927
rect 0 72676 1014 72876
rect 85358 72676 86372 72876
rect 0 71776 1706 72476
rect 84666 71776 86372 72476
rect 0 71376 1014 71576
rect 85358 71376 86372 71576
rect 0 71328 27272 71376
rect 59421 71328 86372 71376
rect 0 71127 86372 71328
rect 0 71076 27272 71127
rect 30403 71126 54622 71127
rect 59421 71076 86372 71127
rect 0 70876 1014 71076
rect 85358 70876 86372 71076
rect 0 69976 1706 70676
rect 84666 69976 86372 70676
rect 0 69576 1014 69776
rect 85358 69576 86372 69776
rect 0 69528 27272 69576
rect 59421 69528 86372 69576
rect 0 69327 86372 69528
rect 0 69276 27272 69327
rect 30403 69326 54622 69327
rect 59421 69276 86372 69327
rect 0 69076 1014 69276
rect 85358 69076 86372 69276
rect 0 68176 1706 68876
rect 84666 68176 86372 68876
rect 0 67776 1014 67976
rect 85358 67776 86372 67976
rect 0 67728 27272 67776
rect 59421 67728 86372 67776
rect 0 67527 86372 67728
rect 0 67476 27272 67527
rect 30403 67526 54622 67527
rect 59421 67476 86372 67527
rect 0 67276 1014 67476
rect 85358 67276 86372 67476
rect 0 66376 1706 67076
rect 84666 66376 86372 67076
rect 0 65976 1014 66176
rect 85358 65976 86372 66176
rect 0 65928 27272 65976
rect 59421 65928 86372 65976
rect 0 65727 86372 65928
rect 0 65676 27272 65727
rect 30403 65726 54622 65727
rect 59421 65676 86372 65727
rect 0 65476 1014 65676
rect 85358 65476 86372 65676
rect 0 64576 1706 65276
rect 84666 64576 86372 65276
rect 0 64176 1014 64376
rect 85358 64176 86372 64376
rect 0 64128 27272 64176
rect 59421 64128 86372 64176
rect 0 63927 86372 64128
rect 0 63876 27272 63927
rect 30403 63926 54622 63927
rect 59421 63876 86372 63927
rect 0 63676 1014 63876
rect 85358 63676 86372 63876
rect 0 62776 1706 63476
rect 84666 62776 86372 63476
rect 0 62376 1014 62576
rect 85358 62376 86372 62576
rect 0 62328 27272 62376
rect 59421 62328 86372 62376
rect 0 62127 86372 62328
rect 0 62076 27272 62127
rect 30403 62126 54622 62127
rect 59421 62076 86372 62127
rect 0 61876 1014 62076
rect 85358 61876 86372 62076
rect 0 60976 1706 61676
rect 84666 60976 86372 61676
rect 0 60576 1014 60776
rect 85358 60576 86372 60776
rect 0 60528 27272 60576
rect 59421 60528 86372 60576
rect 0 60327 86372 60528
rect 0 60276 27272 60327
rect 30403 60326 54622 60327
rect 59421 60276 86372 60327
rect 0 60076 1014 60276
rect 85358 60076 86372 60276
rect 0 59176 1706 59876
rect 84666 59176 86372 59876
rect 0 58776 1014 58976
rect 85358 58776 86372 58976
rect 0 58728 27272 58776
rect 59421 58728 86372 58776
rect 0 58527 86372 58728
rect 0 58476 27272 58527
rect 30403 58526 54622 58527
rect 59421 58476 86372 58527
rect 0 58276 1014 58476
rect 85358 58276 86372 58476
rect 0 57376 1706 58076
rect 84666 57376 86372 58076
rect 0 56976 1014 57176
rect 85358 56976 86372 57176
rect 0 56928 27272 56976
rect 59421 56928 86372 56976
rect 0 56727 86372 56928
rect 0 56676 27272 56727
rect 30403 56726 54622 56727
rect 59421 56676 86372 56727
rect 0 56476 1014 56676
rect 85358 56476 86372 56676
rect 0 55576 1706 56276
rect 84666 55576 86372 56276
rect 0 55176 1014 55376
rect 85358 55176 86372 55376
rect 0 55128 27272 55176
rect 59421 55128 86372 55176
rect 0 54927 86372 55128
rect 0 54876 27272 54927
rect 30403 54926 54622 54927
rect 59421 54876 86372 54927
rect 0 54676 1014 54876
rect 85358 54676 86372 54876
rect 0 53776 1706 54476
rect 84666 53776 86372 54476
rect 0 53376 1014 53576
rect 85358 53376 86372 53576
rect 0 53328 27272 53376
rect 59421 53328 86372 53376
rect 0 53127 86372 53328
rect 0 53076 27272 53127
rect 30403 53126 54622 53127
rect 59421 53076 86372 53127
rect 0 52876 1014 53076
rect 85358 52876 86372 53076
rect 0 51976 1706 52676
rect 84666 51976 86372 52676
rect 0 51576 1014 51776
rect 85358 51576 86372 51776
rect 0 51528 27272 51576
rect 59421 51528 86372 51576
rect 0 51327 86372 51528
rect 0 51276 27272 51327
rect 30403 51326 54622 51327
rect 59421 51276 86372 51327
rect 0 51076 1014 51276
rect 85358 51076 86372 51276
rect 0 50176 1706 50876
rect 84666 50176 86372 50876
rect 0 49776 1014 49976
rect 85358 49776 86372 49976
rect 0 49728 27272 49776
rect 59421 49728 86372 49776
rect 0 49527 86372 49728
rect 0 49476 27272 49527
rect 30403 49526 54622 49527
rect 59421 49476 86372 49527
rect 0 49276 1014 49476
rect 85358 49276 86372 49476
rect 0 48376 1706 49076
rect 84666 48376 86372 49076
rect 0 47976 1014 48176
rect 85358 47976 86372 48176
rect 0 47928 27272 47976
rect 59421 47928 86372 47976
rect 0 47727 86372 47928
rect 0 47676 27272 47727
rect 30403 47726 54622 47727
rect 59421 47676 86372 47727
rect 0 47476 1014 47676
rect 85358 47476 86372 47676
rect 0 46576 1706 47276
rect 84666 46576 86372 47276
rect 0 46176 1014 46376
rect 85358 46176 86372 46376
rect 0 46128 27272 46176
rect 59421 46128 86372 46176
rect 0 45927 86372 46128
rect 0 45876 27272 45927
rect 30403 45926 54622 45927
rect 59421 45876 86372 45927
rect 0 45676 1014 45876
rect 85358 45676 86372 45876
rect 0 44776 1706 45476
rect 84666 44776 86372 45476
rect 0 44376 1014 44576
rect 85358 44376 86372 44576
rect 0 44328 27272 44376
rect 59421 44328 86372 44376
rect 0 44127 86372 44328
rect 0 44076 27272 44127
rect 30403 44126 54622 44127
rect 59421 44076 86372 44127
rect 0 43876 1014 44076
rect 85358 43876 86372 44076
rect 0 42976 1706 43676
rect 84666 42976 86372 43676
rect 0 42576 1014 42776
rect 85358 42576 86372 42776
rect 0 42528 27272 42576
rect 59421 42528 86372 42576
rect 0 42327 86372 42528
rect 0 42276 27272 42327
rect 30403 42326 54622 42327
rect 59421 42276 86372 42327
rect 0 42076 1014 42276
rect 85358 42076 86372 42276
rect 0 41176 1706 41876
rect 84666 41176 86372 41876
rect 0 40776 1014 40976
rect 85358 40776 86372 40976
rect 0 40728 27272 40776
rect 59421 40728 86372 40776
rect 0 40527 86372 40728
rect 0 40476 27272 40527
rect 30403 40526 54622 40527
rect 59421 40476 86372 40527
rect 0 40276 1014 40476
rect 85358 40276 86372 40476
rect 0 39376 1706 40076
rect 84666 39376 86372 40076
rect 0 38976 1014 39176
rect 85358 38976 86372 39176
rect 0 38928 27272 38976
rect 59421 38928 86372 38976
rect 0 38727 86372 38928
rect 0 38676 27272 38727
rect 30403 38726 54622 38727
rect 59421 38676 86372 38727
rect 0 38476 1014 38676
rect 85358 38476 86372 38676
rect 0 37576 1706 38276
rect 84666 37576 86372 38276
rect 0 37176 1014 37376
rect 85358 37176 86372 37376
rect 0 37128 27272 37176
rect 59421 37128 86372 37176
rect 0 36927 86372 37128
rect 0 36876 27272 36927
rect 30403 36926 54622 36927
rect 59421 36876 86372 36927
rect 0 36676 1014 36876
rect 85358 36676 86372 36876
rect 0 35776 1706 36476
rect 84666 35776 86372 36476
rect 0 35126 24917 35326
rect 0 35016 1014 35126
rect 83360 35298 86372 35326
rect 60460 35158 86372 35298
rect 83360 35126 86372 35158
rect 0 34536 27830 35016
rect 85358 35016 86372 35126
rect 58791 34536 86372 35016
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 32318 27214 34124
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 57908 32315 86372 34124
rect 57908 32199 58351 32315
rect 26772 31486 58351 32199
rect 26772 29714 58351 30105
rect 84666 29714 86372 32315
rect 0 29430 86372 29714
rect 0 28412 3011 28416
rect 0 26890 26070 28412
rect 26772 27382 58351 29430
rect 83361 28412 86372 28416
rect 0 26435 27828 26890
rect 6921 26434 8163 26435
rect 17721 26434 18963 26435
rect 23425 26434 27828 26435
rect 58785 26890 86372 28412
rect 57295 26435 86372 26890
rect 66497 26434 67739 26435
rect 77297 26434 78539 26435
rect 0 23380 1706 23938
rect 26770 23380 58348 24278
rect 84666 23380 86372 23938
rect 0 23370 86372 23380
rect 0 22938 27214 23370
rect 27387 22291 57681 23199
rect 57908 22938 86372 23370
rect 57908 22937 83763 22938
rect 27387 22282 27826 22291
rect 0 21827 27826 22282
rect 56078 22282 57681 22291
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 21827 86372 22282
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 19969 86372 20739
rect 0 18016 24250 19969
rect 61807 18016 86372 19969
rect 61825 18015 83763 18016
rect 0 16597 23678 17730
rect 61807 16784 86372 17730
rect 24111 16597 27828 16598
rect 0 15015 27828 16597
rect 46982 15015 86372 16784
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14936 51760 14966
rect 0 14491 47683 14936
rect 0 14329 45977 14491
rect 0 14328 24250 14329
rect 24047 14178 27214 14179
rect 0 13461 27214 14178
rect 0 12846 1706 13461
rect 24047 12934 27214 13461
rect 27387 13760 45977 14329
rect 57295 14328 86372 14968
rect 57295 14327 83763 14328
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 59826 13866 60026 14017
rect 61773 13866 86372 14177
rect 27387 13245 49775 13760
rect 29478 13243 49775 13245
rect 41493 13078 49775 13243
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12570 34761 12846
rect 50228 13461 86372 13866
rect 50228 12846 58421 13461
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12570 86372 12846
rect 0 12046 86372 12570
rect 0 12036 24250 12046
rect 26772 12036 86372 12046
rect 26772 12035 84999 12036
rect 26772 11844 58351 12035
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 10176 27828 11491
rect 29478 11697 58351 11844
rect 29478 10756 41516 11697
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 34741 9972 41516 10756
rect 61825 11491 86372 11493
rect 42261 10740 86372 11491
rect 24047 9515 28729 9516
rect 0 9514 1014 9515
rect 2226 9514 28729 9515
rect 0 8154 28729 9514
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 6982 27828 7595
rect 28178 7652 28729 8154
rect 41857 9502 51430 10420
rect 57295 10176 86372 10740
rect 61805 10175 84482 10176
rect 61825 10173 84482 10175
rect 41857 9165 55482 9502
rect 29513 7900 41397 8582
rect 28178 7084 34622 7652
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 8930 55482 9165
rect 50922 7596 57736 8930
rect 57909 9515 62278 9516
rect 57909 9514 72434 9515
rect 72602 9514 83234 9515
rect 85358 9514 86372 9515
rect 57909 8154 86372 9514
rect 61802 8153 86372 8154
rect 61825 8152 86372 8153
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7392 86372 7595
rect 34860 6984 86372 7392
rect 34860 6592 55482 6984
rect 61802 6982 86372 6984
rect 61802 6981 84787 6982
rect 61825 6980 84787 6981
rect 34860 6573 41397 6592
rect 29458 6199 41397 6573
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 0 5766 34622 6177
rect 23687 5629 27214 5630
rect 0 5175 27214 5629
rect 29458 5665 34622 5766
rect 50922 6199 55482 6592
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 50922 5766 86372 6198
rect 50922 5605 55482 5766
rect 0 5174 24250 5175
rect 0 5173 3011 5174
rect 0 4515 1712 5173
rect 57909 5629 62429 5630
rect 57909 5175 86372 5629
rect 61802 5174 86372 5175
rect 83361 5173 86372 5174
rect 57909 4619 62429 4621
rect 23909 4515 62429 4619
rect 84660 4515 86372 5173
rect 0 4166 86372 4515
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 61788 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3772 61215 3875
rect 0 3524 86372 3772
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 0 2854 1014 3420
rect 60886 3420 86372 3524
rect 85358 2854 86372 3420
rect 0 2502 86372 2854
rect 0 1232 86372 2232
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
<< obsm3 >>
rect 0 96232 1345 96976
rect 2457 96312 2570 96976
rect 3682 96312 4081 96976
rect 2457 96232 4081 96312
rect 5193 96312 5306 96976
rect 6418 96312 6745 96976
rect 5193 96232 6745 96312
rect 7857 96312 7970 96976
rect 9082 96312 9481 96976
rect 7857 96232 9481 96312
rect 10593 96312 10706 96976
rect 11818 96312 12145 96976
rect 10593 96232 12145 96312
rect 13257 96312 13370 96976
rect 14482 96312 14881 96976
rect 13257 96232 14881 96312
rect 15993 96312 16106 96976
rect 17218 96312 17545 96976
rect 15993 96232 17545 96312
rect 18657 96312 18770 96976
rect 19882 96312 20597 96976
rect 18657 96232 20597 96312
rect 21709 96312 22202 96976
rect 23314 96312 23427 96976
rect 21709 96232 23427 96312
rect 24539 96312 25102 96976
rect 26214 96312 26516 96976
rect 24539 96232 26516 96312
rect 27628 96312 27821 96976
rect 28933 96312 29217 96976
rect 30329 96312 30654 96976
rect 27628 96232 30654 96312
rect 31766 96312 32325 96976
rect 33437 96312 33968 96976
rect 35080 96312 35359 96976
rect 31766 96232 35359 96312
rect 36471 96312 36892 96976
rect 38004 96312 38529 96976
rect 36471 96232 38529 96312
rect 39641 96312 39826 96976
rect 40938 96312 41174 96976
rect 39641 96232 41174 96312
rect 42286 96312 42374 96976
rect 43486 96312 43657 96976
rect 44769 96312 45013 96976
rect 42286 96232 45013 96312
rect 46125 96232 46257 96976
rect 47369 96312 47482 96976
rect 48594 96312 48845 96976
rect 47369 96232 48845 96312
rect 49957 96312 50409 96976
rect 51521 96312 52513 96976
rect 49957 96232 52513 96312
rect 53625 96232 54206 96976
rect 55318 96312 55934 96976
rect 57046 96312 57491 96976
rect 55318 96232 57491 96312
rect 58603 96312 58735 96976
rect 59847 96312 60921 96976
rect 58603 96232 60921 96312
rect 62033 96312 62146 96976
rect 63258 96312 63657 96976
rect 62033 96232 63657 96312
rect 64769 96312 64882 96976
rect 65994 96312 66321 96976
rect 64769 96232 66321 96312
rect 67433 96312 67546 96976
rect 68658 96312 69057 96976
rect 67433 96232 69057 96312
rect 70169 96312 70282 96976
rect 71394 96312 71721 96976
rect 70169 96232 71721 96312
rect 72833 96312 72946 96976
rect 74058 96312 74457 96976
rect 72833 96232 74457 96312
rect 75569 96312 75682 96976
rect 76794 96312 77121 96976
rect 75569 96232 77121 96312
rect 78233 96312 78346 96976
rect 79458 96312 80173 96976
rect 78233 96232 80173 96312
rect 81285 96312 81778 96976
rect 82890 96312 83003 96976
rect 81285 96232 83003 96312
rect 84115 96232 84610 96976
rect 85722 96232 86372 96976
rect 0 95032 86372 95120
rect 1070 94841 85302 95032
rect 1070 94832 25320 94841
rect 26004 94832 58799 94841
rect 59483 94832 85302 94841
rect 27328 94784 58799 94832
rect 27328 94470 30346 94471
rect 54678 94470 58799 94471
rect 27328 94420 58799 94470
rect 1070 94405 25320 94420
rect 26004 94405 58799 94420
rect 59483 94405 85302 94420
rect 1070 94220 85302 94405
rect 0 94132 86372 94220
rect 1762 93320 84610 94132
rect 0 93232 86372 93320
rect 1070 93032 85302 93232
rect 27328 92984 59365 93032
rect 27328 92670 30347 92671
rect 54678 92670 59365 92671
rect 27328 92620 59365 92670
rect 1070 92420 85302 92620
rect 0 92332 86372 92420
rect 1762 91520 84610 92332
rect 0 91432 86372 91520
rect 1070 91232 85302 91432
rect 27328 91184 59365 91232
rect 27328 90870 30347 90871
rect 54678 90870 59365 90871
rect 27328 90820 59365 90870
rect 1070 90620 85302 90820
rect 0 90532 86372 90620
rect 1762 89720 84610 90532
rect 0 89632 86372 89720
rect 1070 89432 85302 89632
rect 27328 89384 59365 89432
rect 27328 89070 30347 89071
rect 54678 89070 59365 89071
rect 27328 89020 59365 89070
rect 1070 88820 85302 89020
rect 0 88732 86372 88820
rect 1762 87920 84610 88732
rect 0 87832 86372 87920
rect 1070 87632 85302 87832
rect 27328 87584 59365 87632
rect 27328 87270 30347 87271
rect 54678 87270 59365 87271
rect 27328 87220 59365 87270
rect 1070 87020 85302 87220
rect 0 86932 86372 87020
rect 1762 86120 84610 86932
rect 0 86032 86372 86120
rect 1070 85832 85302 86032
rect 27328 85784 59365 85832
rect 27328 85470 30347 85471
rect 54678 85470 59365 85471
rect 27328 85420 59365 85470
rect 1070 85220 85302 85420
rect 0 85132 86372 85220
rect 1762 84320 84610 85132
rect 0 84232 86372 84320
rect 1070 84032 85302 84232
rect 27328 83984 59365 84032
rect 27328 83670 30347 83671
rect 54678 83670 59365 83671
rect 27328 83620 59365 83670
rect 1070 83420 85302 83620
rect 0 83332 86372 83420
rect 1762 82520 84610 83332
rect 0 82432 86372 82520
rect 1070 82232 85302 82432
rect 27328 82184 59365 82232
rect 27328 81870 30347 81871
rect 54678 81870 59365 81871
rect 27328 81820 59365 81870
rect 1070 81620 85302 81820
rect 0 81532 86372 81620
rect 1762 80720 84610 81532
rect 0 80632 86372 80720
rect 1070 80432 85302 80632
rect 27328 80384 59365 80432
rect 27328 80070 30347 80071
rect 54678 80070 59365 80071
rect 27328 80020 59365 80070
rect 1070 79820 85302 80020
rect 0 79732 86372 79820
rect 1762 78920 84610 79732
rect 0 78832 86372 78920
rect 1070 78632 85302 78832
rect 27328 78584 59365 78632
rect 27328 78270 30347 78271
rect 54678 78270 59365 78271
rect 27328 78220 59365 78270
rect 1070 78020 85302 78220
rect 0 77932 86372 78020
rect 1762 77120 84610 77932
rect 0 77032 86372 77120
rect 1070 76832 85302 77032
rect 27328 76784 59365 76832
rect 27328 76470 30347 76471
rect 54678 76470 59365 76471
rect 27328 76420 59365 76470
rect 1070 76220 85302 76420
rect 0 76132 86372 76220
rect 1762 75320 84610 76132
rect 0 75232 86372 75320
rect 1070 75032 85302 75232
rect 27328 74984 59365 75032
rect 27328 74670 30347 74671
rect 54678 74670 59365 74671
rect 27328 74620 59365 74670
rect 1070 74420 85302 74620
rect 0 74332 86372 74420
rect 1762 73520 84610 74332
rect 0 73432 86372 73520
rect 1070 73232 85302 73432
rect 27328 73184 59365 73232
rect 27328 72870 30347 72871
rect 54678 72870 59365 72871
rect 27328 72820 59365 72870
rect 1070 72620 85302 72820
rect 0 72532 86372 72620
rect 1762 71720 84610 72532
rect 0 71632 86372 71720
rect 1070 71432 85302 71632
rect 27328 71384 59365 71432
rect 27328 71070 30347 71071
rect 54678 71070 59365 71071
rect 27328 71020 59365 71070
rect 1070 70820 85302 71020
rect 0 70732 86372 70820
rect 1762 69920 84610 70732
rect 0 69832 86372 69920
rect 1070 69632 85302 69832
rect 27328 69584 59365 69632
rect 27328 69270 30347 69271
rect 54678 69270 59365 69271
rect 27328 69220 59365 69270
rect 1070 69020 85302 69220
rect 0 68932 86372 69020
rect 1762 68120 84610 68932
rect 0 68032 86372 68120
rect 1070 67832 85302 68032
rect 27328 67784 59365 67832
rect 27328 67470 30347 67471
rect 54678 67470 59365 67471
rect 27328 67420 59365 67470
rect 1070 67220 85302 67420
rect 0 67132 86372 67220
rect 1762 66320 84610 67132
rect 0 66232 86372 66320
rect 1070 66032 85302 66232
rect 27328 65984 59365 66032
rect 27328 65670 30347 65671
rect 54678 65670 59365 65671
rect 27328 65620 59365 65670
rect 1070 65420 85302 65620
rect 0 65332 86372 65420
rect 1762 64520 84610 65332
rect 0 64432 86372 64520
rect 1070 64232 85302 64432
rect 27328 64184 59365 64232
rect 27328 63870 30347 63871
rect 54678 63870 59365 63871
rect 27328 63820 59365 63870
rect 1070 63620 85302 63820
rect 0 63532 86372 63620
rect 1762 62720 84610 63532
rect 0 62632 86372 62720
rect 1070 62432 85302 62632
rect 27328 62384 59365 62432
rect 27328 62070 30347 62071
rect 54678 62070 59365 62071
rect 27328 62020 59365 62070
rect 1070 61820 85302 62020
rect 0 61732 86372 61820
rect 1762 60920 84610 61732
rect 0 60832 86372 60920
rect 1070 60632 85302 60832
rect 27328 60584 59365 60632
rect 27328 60270 30347 60271
rect 54678 60270 59365 60271
rect 27328 60220 59365 60270
rect 1070 60020 85302 60220
rect 0 59932 86372 60020
rect 1762 59120 84610 59932
rect 0 59032 86372 59120
rect 1070 58832 85302 59032
rect 27328 58784 59365 58832
rect 27328 58470 30347 58471
rect 54678 58470 59365 58471
rect 27328 58420 59365 58470
rect 1070 58220 85302 58420
rect 0 58132 86372 58220
rect 1762 57320 84610 58132
rect 0 57232 86372 57320
rect 1070 57032 85302 57232
rect 27328 56984 59365 57032
rect 27328 56670 30347 56671
rect 54678 56670 59365 56671
rect 27328 56620 59365 56670
rect 1070 56420 85302 56620
rect 0 56332 86372 56420
rect 1762 55520 84610 56332
rect 0 55432 86372 55520
rect 1070 55232 85302 55432
rect 27328 55184 59365 55232
rect 27328 54870 30347 54871
rect 54678 54870 59365 54871
rect 27328 54820 59365 54870
rect 1070 54620 85302 54820
rect 0 54532 86372 54620
rect 1762 53720 84610 54532
rect 0 53632 86372 53720
rect 1070 53432 85302 53632
rect 27328 53384 59365 53432
rect 27328 53070 30347 53071
rect 54678 53070 59365 53071
rect 27328 53020 59365 53070
rect 1070 52820 85302 53020
rect 0 52732 86372 52820
rect 1762 51920 84610 52732
rect 0 51832 86372 51920
rect 1070 51632 85302 51832
rect 27328 51584 59365 51632
rect 27328 51270 30347 51271
rect 54678 51270 59365 51271
rect 27328 51220 59365 51270
rect 1070 51020 85302 51220
rect 0 50932 86372 51020
rect 1762 50120 84610 50932
rect 0 50032 86372 50120
rect 1070 49832 85302 50032
rect 27328 49784 59365 49832
rect 27328 49470 30347 49471
rect 54678 49470 59365 49471
rect 27328 49420 59365 49470
rect 1070 49220 85302 49420
rect 0 49132 86372 49220
rect 1762 48320 84610 49132
rect 0 48232 86372 48320
rect 1070 48032 85302 48232
rect 27328 47984 59365 48032
rect 27328 47670 30347 47671
rect 54678 47670 59365 47671
rect 27328 47620 59365 47670
rect 1070 47420 85302 47620
rect 0 47332 86372 47420
rect 1762 46520 84610 47332
rect 0 46432 86372 46520
rect 1070 46232 85302 46432
rect 27328 46184 59365 46232
rect 27328 45870 30347 45871
rect 54678 45870 59365 45871
rect 27328 45820 59365 45870
rect 1070 45620 85302 45820
rect 0 45532 86372 45620
rect 1762 44720 84610 45532
rect 0 44632 86372 44720
rect 1070 44432 85302 44632
rect 27328 44384 59365 44432
rect 27328 44070 30347 44071
rect 54678 44070 59365 44071
rect 27328 44020 59365 44070
rect 1070 43820 85302 44020
rect 0 43732 86372 43820
rect 1762 42920 84610 43732
rect 0 42832 86372 42920
rect 1070 42632 85302 42832
rect 27328 42584 59365 42632
rect 27328 42270 30347 42271
rect 54678 42270 59365 42271
rect 27328 42220 59365 42270
rect 1070 42020 85302 42220
rect 0 41932 86372 42020
rect 1762 41120 84610 41932
rect 0 41032 86372 41120
rect 1070 40832 85302 41032
rect 27328 40784 59365 40832
rect 27328 40470 30347 40471
rect 54678 40470 59365 40471
rect 27328 40420 59365 40470
rect 1070 40220 85302 40420
rect 0 40132 86372 40220
rect 1762 39320 84610 40132
rect 0 39232 86372 39320
rect 1070 39032 85302 39232
rect 27328 38984 59365 39032
rect 27328 38670 30347 38671
rect 54678 38670 59365 38671
rect 27328 38620 59365 38670
rect 1070 38420 85302 38620
rect 0 38332 86372 38420
rect 1762 37520 84610 38332
rect 0 37432 86372 37520
rect 1070 37232 85302 37432
rect 27328 37184 59365 37232
rect 27328 36870 30347 36871
rect 54678 36870 59365 36871
rect 27328 36820 59365 36870
rect 1070 36620 85302 36820
rect 0 36532 86372 36620
rect 1762 35720 84610 36532
rect 0 35382 86372 35720
rect 24973 35354 83304 35382
rect 24973 35102 60404 35354
rect 24973 35072 83304 35102
rect 27886 34480 58735 35072
rect 0 34182 86372 34480
rect 0 34181 2039 34182
rect 2244 34181 86372 34182
rect 25141 34180 61797 34181
rect 72439 34180 72597 34181
rect 27270 32262 57852 34180
rect 25141 32260 57852 32262
rect 3067 32259 57852 32260
rect 1762 32255 57852 32259
rect 1762 31430 26716 32255
rect 58407 31430 84610 32259
rect 1762 30161 84610 31430
rect 1762 29770 26716 30161
rect 58407 29770 84610 30161
rect 0 28472 26716 29374
rect 3067 28468 26716 28472
rect 26126 27326 26716 28468
rect 58407 28472 86372 29374
rect 58407 28468 83305 28472
rect 58407 27326 58729 28468
rect 26126 26946 58729 27326
rect 27884 26379 57239 26946
rect 0 26378 6865 26379
rect 8219 26378 17665 26379
rect 19019 26378 23369 26379
rect 27884 26378 66441 26379
rect 67795 26378 77241 26379
rect 78595 26378 86372 26379
rect 0 24334 86372 26378
rect 0 23994 26714 24334
rect 1762 23436 26714 23994
rect 58404 23994 86372 24334
rect 58404 23436 84610 23994
rect 27270 23255 57852 23314
rect 27270 22882 27331 23255
rect 0 22338 27331 22882
rect 57737 22881 57852 23255
rect 83819 22881 86372 22882
rect 57737 22338 86372 22881
rect 1070 21770 23980 21771
rect 27882 21770 56022 22235
rect 83819 21770 85302 21771
rect 1070 21764 85302 21770
rect 1070 21763 44376 21764
rect 1070 21681 29465 21763
rect 1070 21226 29457 21681
rect 0 20795 29457 21226
rect 55701 21226 85302 21764
rect 55701 20795 86372 21226
rect 24306 17960 61751 19913
rect 0 17959 61769 17960
rect 83819 17959 86372 17960
rect 0 17786 86372 17959
rect 23734 16840 61751 17786
rect 23734 16654 46926 16840
rect 23734 16653 24055 16654
rect 27884 15071 46926 16654
rect 55701 14910 57239 14912
rect 51816 14880 57239 14910
rect 47739 14435 57239 14880
rect 24306 14272 27331 14273
rect 0 14235 27331 14272
rect 0 14234 23991 14235
rect 1762 12903 23991 13405
rect 27270 13189 27331 14235
rect 46033 14271 57239 14435
rect 83819 14271 86372 14272
rect 46033 14235 86372 14271
rect 46033 14234 83113 14235
rect 84277 14234 86372 14235
rect 46033 14233 61751 14234
rect 72485 14233 72551 14234
rect 46033 14073 61717 14233
rect 46033 13922 59770 14073
rect 46033 13816 50172 13922
rect 60082 13922 61717 14073
rect 27270 13187 29422 13189
rect 27270 13022 41437 13187
rect 49831 13022 50172 13816
rect 27270 12990 50172 13022
rect 1762 12902 23765 12903
rect 34817 12626 50172 12990
rect 58477 12902 59770 13405
rect 60082 12903 84610 13405
rect 60082 12902 83113 12903
rect 84277 12902 84610 12903
rect 24306 11980 26716 11990
rect 0 11788 26716 11980
rect 85055 11979 86372 11980
rect 0 11549 29422 11788
rect 3067 11547 23991 11549
rect 27884 10700 29422 11549
rect 58407 11641 86372 11979
rect 27884 10120 34685 10700
rect 0 10119 2173 10120
rect 0 10118 2193 10119
rect 24306 10118 34685 10120
rect 0 9916 34685 10118
rect 41572 11549 86372 11641
rect 41572 11547 61769 11549
rect 41572 10684 42205 11547
rect 41572 10476 57239 10684
rect 41572 9916 41801 10476
rect 0 9572 41801 9916
rect 0 9571 23991 9572
rect 1070 9570 2170 9571
rect 24306 8097 28122 8098
rect 3067 8096 28122 8097
rect 0 7652 28122 8096
rect 3067 7651 23569 7652
rect 27884 7028 28122 7652
rect 28785 9109 41801 9572
rect 51486 10120 57239 10476
rect 51486 10119 61749 10120
rect 51486 10117 61769 10119
rect 84538 10117 86372 10120
rect 51486 9572 86372 10117
rect 51486 9558 57853 9572
rect 62334 9571 86372 9572
rect 72490 9570 72546 9571
rect 83290 9570 85302 9571
rect 28785 8638 50866 9109
rect 28785 7844 29457 8638
rect 28785 7708 34804 7844
rect 27884 6926 29481 7028
rect 1070 6925 2170 6926
rect 1070 6924 2193 6925
rect 24306 6924 29481 6926
rect 1070 6688 29481 6924
rect 34678 6688 34804 7708
rect 1070 6629 34804 6688
rect 41453 7448 50866 8638
rect 55538 8986 57853 9558
rect 57792 8098 57853 8986
rect 57792 8097 61746 8098
rect 57792 8096 61769 8097
rect 57792 7652 86372 8096
rect 62803 7651 83305 7652
rect 1070 6255 29402 6629
rect 3067 6254 23631 6255
rect 41453 6121 50866 6536
rect 0 5686 29402 5710
rect 0 5685 23631 5686
rect 27270 5609 29402 5686
rect 34678 5609 50866 6121
rect 27270 5549 50866 5609
rect 55538 6925 61746 6928
rect 55538 6924 61769 6925
rect 84843 6924 85302 6926
rect 55538 6255 85302 6924
rect 62485 6254 83305 6255
rect 55538 5686 86372 5710
rect 55538 5549 57853 5686
rect 62485 5685 86372 5686
rect 27270 5119 57853 5549
rect 24306 5118 61746 5119
rect 3067 5117 83305 5118
rect 1768 4677 84604 5117
rect 1768 4675 57853 4677
rect 1768 4571 23853 4675
rect 62485 4571 84604 4677
rect 59379 4108 61732 4110
rect 24397 4004 61732 4108
rect 0 3932 86372 4004
rect 0 3931 27382 3932
rect 27834 3931 28708 3932
rect 28950 3931 41718 3932
rect 41960 3931 42243 3932
rect 42485 3931 46817 3932
rect 47059 3931 47265 3932
rect 47507 3931 47713 3932
rect 47955 3931 48161 3932
rect 48403 3931 57289 3932
rect 0 3828 23853 3931
rect 61271 3828 86372 3932
rect 24397 3365 60830 3468
rect 3067 3364 60830 3365
rect 1070 2910 85302 3364
rect 0 2288 86372 2446
rect 0 0 650 1176
rect 1762 0 1983 1176
rect 3095 0 3386 1176
rect 4498 988 5786 1176
rect 4498 0 4586 988
rect 5698 0 5786 988
rect 6898 0 6986 1176
rect 8098 0 8186 1176
rect 9298 988 10586 1176
rect 9298 0 9386 988
rect 10498 0 10586 988
rect 11698 0 12387 1176
rect 13499 0 14186 1176
rect 15298 988 16586 1176
rect 15298 0 15386 988
rect 16498 0 16586 988
rect 17698 0 17786 1176
rect 18898 0 18986 1176
rect 20098 988 21854 1176
rect 20098 0 20186 988
rect 21298 0 21854 988
rect 22966 0 23054 1176
rect 24166 0 24354 1176
rect 25466 0 25654 1176
rect 26766 0 26954 1176
rect 28066 0 28254 1176
rect 29366 0 29554 1176
rect 30666 988 35975 1176
rect 30666 0 31268 988
rect 32380 0 32966 988
rect 34078 0 34775 988
rect 35887 0 35975 988
rect 37087 988 39172 1176
rect 37087 0 37972 988
rect 39084 0 39172 988
rect 40284 988 42377 1176
rect 40284 0 41177 988
rect 42289 0 42377 988
rect 43489 988 44777 1176
rect 43489 0 43577 988
rect 44689 0 44777 988
rect 45889 988 47177 1176
rect 45889 0 45977 988
rect 47089 0 47177 988
rect 48289 0 48510 1176
rect 49622 0 49820 1176
rect 50932 988 54402 1176
rect 50932 0 51177 988
rect 52289 0 52422 988
rect 53534 0 54402 988
rect 55514 0 55702 1176
rect 56814 0 57002 1176
rect 58114 0 58302 1176
rect 59414 0 59602 1176
rect 60714 0 60902 1176
rect 62014 0 62239 1176
rect 63351 988 65362 1176
rect 63351 0 64162 988
rect 65274 0 65362 988
rect 66474 0 66562 1176
rect 67674 0 67762 1176
rect 68874 988 70162 1176
rect 68874 0 68962 988
rect 70074 0 70162 988
rect 71274 0 71961 1176
rect 73073 0 73762 1176
rect 74874 988 76162 1176
rect 74874 0 74962 988
rect 76074 0 76162 988
rect 77274 0 77362 1176
rect 78474 0 78562 1176
rect 79674 988 80962 1176
rect 79674 0 79762 988
rect 80874 0 80962 988
rect 82074 0 82363 1176
rect 83475 0 84610 1176
rect 85722 0 86372 1176
<< labels >>
rlabel metal2 s 34243 0 34467 200 6 A[0]
port 9 nsew signal input
rlabel metal2 s 32552 0 32776 200 6 A[1]
port 8 nsew signal input
rlabel metal2 s 30859 0 31083 200 6 A[2]
port 7 nsew signal input
rlabel metal2 s 56265 0 56489 200 6 A[3]
port 6 nsew signal input
rlabel metal2 s 55164 0 55388 200 6 A[4]
port 5 nsew signal input
rlabel metal2 s 54417 0 54641 200 6 A[5]
port 4 nsew signal input
rlabel metal2 s 53772 0 53996 200 6 A[6]
port 3 nsew signal input
rlabel metal2 s 29705 0 29929 200 6 A[7]
port 2 nsew signal input
rlabel metal2 s 29006 0 29230 200 6 A[8]
port 1 nsew signal input
rlabel metal2 s 50342 0 50566 200 6 CEN
port 10 nsew signal input
rlabel metal2 s 27936 0 28160 200 6 CLK
port 11 nsew signal input
rlabel metal2 s 1864 0 2088 200 6 D[0]
port 19 nsew signal input
rlabel metal2 s 12206 0 12430 200 6 D[1]
port 18 nsew signal input
rlabel metal2 s 13454 0 13678 200 6 D[2]
port 17 nsew signal input
rlabel metal2 s 23795 0 24019 200 6 D[3]
port 16 nsew signal input
rlabel metal2 s 61447 0 61671 200 6 D[4]
port 15 nsew signal input
rlabel metal2 s 71782 0 72006 200 6 D[5]
port 14 nsew signal input
rlabel metal2 s 73030 0 73254 200 6 D[6]
port 13 nsew signal input
rlabel metal2 s 83372 0 83596 200 6 D[7]
port 12 nsew signal input
rlabel metal2 s 40588 0 40812 200 6 GWEN
port 20 nsew signal input
rlabel metal2 s 3380 0 3604 200 6 Q[0]
port 28 nsew signal output
rlabel metal2 s 11533 0 11757 200 6 Q[1]
port 27 nsew signal output
rlabel metal2 s 14127 0 14351 200 6 Q[2]
port 26 nsew signal output
rlabel metal2 s 22279 0 22503 200 6 Q[3]
port 25 nsew signal output
rlabel metal2 s 62958 0 63182 200 6 Q[4]
port 24 nsew signal output
rlabel metal2 s 71109 0 71333 200 6 Q[5]
port 23 nsew signal output
rlabel metal2 s 73703 0 73927 200 6 Q[6]
port 22 nsew signal output
rlabel metal2 s 81855 0 82079 200 6 Q[7]
port 21 nsew signal output
rlabel metal2 s 2539 0 2763 200 6 WEN[0]
port 38 nsew signal input
rlabel metal2 s 12604 0 12828 200 6 WEN[1]
port 37 nsew signal input
rlabel metal2 s 13054 0 13278 200 6 WEN[2]
port 36 nsew signal input
rlabel metal2 s 23404 0 23628 200 6 WEN[3]
port 35 nsew signal input
rlabel metal2 s 62115 0 62339 200 6 WEN[4]
port 34 nsew signal input
rlabel metal2 s 72180 0 72404 200 6 WEN[5]
port 33 nsew signal input
rlabel metal2 s 72630 0 72854 200 6 WEN[6]
port 32 nsew signal input
rlabel metal2 s 82695 0 82919 200 6 WEN[7]
port 31 nsew signal input
rlabel metal3 s 0 93376 1706 94076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 91576 1706 92276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 89776 1706 90476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 87976 1706 88676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 86176 1706 86876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 84376 1706 85076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 82576 1706 83276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 80776 1706 81476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 78976 1706 79676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 77176 1706 77876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 75376 1706 76076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 73576 1706 74276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 71776 1706 72476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 69976 1706 70676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 68176 1706 68876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 66376 1706 67076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 64576 1706 65276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 62776 1706 63476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 60976 1706 61676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 59176 1706 59876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 57376 1706 58076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 55576 1706 56276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 53776 1706 54476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 51976 1706 52676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 50176 1706 50876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 48376 1706 49076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 46576 1706 47276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 44776 1706 45476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 42976 1706 43676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 41176 1706 41876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 39376 1706 40076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 37576 1706 38276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 35776 1706 36476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 8152 1014 9515 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 8152 3011 9514 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 2226 8154 28729 9515 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 8153 24250 9514 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 28178 7084 28729 9516 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 24047 8154 28729 9516 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 29537 6744 34622 7652 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 28178 7084 34622 7652 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 1401 95176 2401 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 4137 95176 5137 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 6801 95176 7801 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 9537 95176 10537 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 12201 95176 13201 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 14937 95176 15937 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 17601 95176 18601 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 20653 95176 21653 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23483 95176 24483 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 26572 95176 27572 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 30710 95176 31710 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 35415 95176 36415 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 38585 95176 39585 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 41230 95176 42230 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 45069 95176 46069 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 46313 95176 47313 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 48901 95176 49901 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 52569 95176 53569 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 54262 95176 55262 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57547 95176 58547 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 60977 95176 61977 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 63713 95176 64713 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 66377 95176 67377 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 69113 95176 70113 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 71777 95176 72777 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 74513 95176 75513 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 77177 95176 78177 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 80229 95176 81229 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 83059 95176 84059 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 95176 85666 96976 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 95176 86372 96176 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 93376 86372 94076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 91576 86372 92276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 89776 86372 90476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 87976 86372 88676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 86176 86372 86876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 84376 86372 85076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 82576 86372 83276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 80776 86372 81476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 78976 86372 79676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 77176 86372 77876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 75376 86372 76076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 73576 86372 74276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 71776 86372 72476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 69976 86372 70676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 68176 86372 68876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 66376 86372 67076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 64576 86372 65276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 62776 86372 63476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 60976 86372 61676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 59176 86372 59876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 57376 86372 58076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 55576 86372 56276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 53776 86372 54476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 51976 86372 52676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 50176 86372 50876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 48376 86372 49076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 46576 86372 47276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 44776 86372 45476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 42976 86372 43676 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 41176 86372 41876 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 39376 86372 40076 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 37576 86372 38276 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 35776 86372 36476 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 29430 1706 34125 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 2095 32315 2188 34126 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 32315 3011 34125 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 32316 25085 34125 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 32318 27214 34124 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 26772 31486 58351 32199 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 26772 27382 58351 30105 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57908 31486 58351 34124 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61853 32315 72383 34125 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57908 32315 86372 34124 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 29430 86372 29714 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 29430 86372 34125 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 72653 32315 86372 34125 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 22938 1706 23938 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 22938 27214 23380 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 26770 23370 58348 24278 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57908 22937 83763 23380 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57908 22938 86372 23380 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 22938 86372 23938 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 18016 24250 20739 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 29513 19969 55645 21625 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 29521 19969 55645 21707 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 44432 19969 55645 21708 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61825 18015 83763 20739 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61807 18016 86372 20739 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 19969 86372 20739 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 12036 1706 14178 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23821 12046 34761 12847 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 13461 27214 14178 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 12036 24250 12846 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 24047 12046 27214 14179 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 24047 12046 34761 12934 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 34741 9972 41516 12570 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 29478 10756 41516 12570 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 29478 11697 58351 12570 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 26772 11844 58351 12570 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 50228 12035 58421 13866 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 59826 12035 60026 14017 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 50228 13461 86372 13866 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61807 13461 72429 14178 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61773 13461 86372 14177 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 83169 12035 84221 12847 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 83169 13461 84221 14179 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 50228 12036 86372 12846 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 26772 12035 84999 12570 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 12036 86372 14178 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 72607 13461 86372 14178 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61802 8153 86372 9514 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57909 8154 62278 9516 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57909 8154 72434 9515 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 72602 8152 83234 9515 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61825 8152 86372 9514 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 85358 8152 86372 9515 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 4060 1712 5629 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 5173 3011 5629 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 5174 24250 5629 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 4060 24341 4515 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23687 5175 27214 5630 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61788 4060 86372 4515 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61802 5174 86372 5629 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 6 VDD
port 29 nsew power bidirectional
rlabel metal3 s 2626 96368 3626 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 4642 0 5642 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 5362 96368 6362 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 8026 96368 9026 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 9442 0 10442 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 10762 96368 11762 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 13426 96368 14426 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 15442 0 16442 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 16162 96368 17162 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 18826 96368 19826 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 20242 0 21242 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 22258 96368 23258 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 25158 96368 26158 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 26435 3011 28416 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 6921 26434 8163 28412 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 17721 26434 18963 28412 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 26435 26070 28412 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23425 26434 27828 26890 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 10176 3011 11493 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 2249 10174 24250 11491 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 2229 10175 24250 11491 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 24047 10176 27828 11493 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 34536 1014 35326 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 35126 24917 35326 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 34536 27830 35016 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27877 96368 28877 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29273 96368 30273 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 31324 0 32324 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 32381 96368 33381 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 33022 0 34022 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 34024 96368 35024 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 34831 0 35831 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 36948 96368 37948 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 38028 0 39028 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 39882 96368 40882 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41233 0 42233 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 42430 96368 43430 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 43633 0 44633 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 43713 96368 44713 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 46033 0 47033 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 47538 96368 48538 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50465 96368 51465 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 51233 0 52233 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 52478 0 53478 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 55990 96368 56990 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58791 96368 59791 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 62202 96368 63202 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 64218 0 65218 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 64938 96368 65938 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 67602 96368 68602 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 69018 0 70018 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 70338 96368 71338 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 73002 96368 74002 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 75018 0 76018 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 75738 96368 76738 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 78402 96368 79402 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 79818 0 80818 932 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 81834 96368 82834 96976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 94276 1014 94976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 25376 94461 25948 94785 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 94476 27272 94776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30402 94526 54622 94728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 94527 86372 94728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58855 94461 59427 94785 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58855 94476 86372 94776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 94276 86372 94976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 92476 1014 93176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 92676 27272 92976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 92726 54622 92928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 92727 86372 92928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 92676 86372 92976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 92476 86372 93176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 90676 1014 91376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 90876 27272 91176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 90926 54622 91128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 90927 86372 91128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 90876 86372 91176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 90676 86372 91376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 88876 1014 89576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 89076 27272 89376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 89126 54622 89328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 89127 86372 89328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 89076 86372 89376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 88876 86372 89576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 87076 1014 87776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 87276 27272 87576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 87326 54622 87528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 87327 86372 87528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 87276 86372 87576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 87076 86372 87776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 85276 1014 85976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 85476 27272 85776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 85526 54622 85728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 85527 86372 85728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 85476 86372 85776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 85276 86372 85976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 83476 1014 84176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 83676 27272 83976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 83726 54622 83928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 83727 86372 83928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 83676 86372 83976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 83476 86372 84176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 81676 1014 82376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 81876 27272 82176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 81926 54622 82128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 81927 86372 82128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 81876 86372 82176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 81676 86372 82376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 79876 1014 80576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 80076 27272 80376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 80126 54622 80328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 80127 86372 80328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 80076 86372 80376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 79876 86372 80576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 78076 1014 78776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 78276 27272 78576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 78326 54622 78528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 78327 86372 78528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 78276 86372 78576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 78076 86372 78776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 76276 1014 76976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 76476 27272 76776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 76526 54622 76728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 76527 86372 76728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 76476 86372 76776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 76276 86372 76976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 74476 1014 75176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 74676 27272 74976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 74726 54622 74928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 74727 86372 74928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 74676 86372 74976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 74476 86372 75176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72676 1014 73376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72876 27272 73176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 72926 54622 73128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72927 86372 73128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 72876 86372 73176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 72676 86372 73376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 70876 1014 71576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 71076 27272 71376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 71126 54622 71328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 71127 86372 71328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 71076 86372 71376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 70876 86372 71576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69076 1014 69776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69276 27272 69576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 69326 54622 69528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69327 86372 69528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 69276 86372 69576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 69076 86372 69776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67276 1014 67976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67476 27272 67776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 67526 54622 67728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67527 86372 67728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 67476 86372 67776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 67276 86372 67976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65476 1014 66176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65676 27272 65976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 65726 54622 65928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65727 86372 65928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 65676 86372 65976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 65476 86372 66176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63676 1014 64376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63876 27272 64176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 63926 54622 64128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63927 86372 64128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 63876 86372 64176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 63676 86372 64376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 61876 1014 62576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 62076 27272 62376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 62126 54622 62328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 62127 86372 62328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 62076 86372 62376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 61876 86372 62576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60076 1014 60776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60276 27272 60576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 60326 54622 60528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60327 86372 60528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 60276 86372 60576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 60076 86372 60776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58276 1014 58976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58476 27272 58776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 58526 54622 58728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58527 86372 58728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 58476 86372 58776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 58276 86372 58976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56476 1014 57176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56676 27272 56976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 56726 54622 56928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56727 86372 56928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 56676 86372 56976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 56476 86372 57176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54676 1014 55376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54876 27272 55176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 54926 54622 55128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54927 86372 55128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 54876 86372 55176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 54676 86372 55376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 52876 1014 53576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 53076 27272 53376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 53126 54622 53328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 53127 86372 53328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 53076 86372 53376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 52876 86372 53576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51076 1014 51776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51276 27272 51576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 51326 54622 51528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51327 86372 51528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 51276 86372 51576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 51076 86372 51776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49276 1014 49976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49476 27272 49776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 49526 54622 49728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49527 86372 49728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 49476 86372 49776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 49276 86372 49976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47476 1014 48176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47676 27272 47976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 47726 54622 47928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47727 86372 47928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 47676 86372 47976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 47476 86372 48176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45676 1014 46376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45876 27272 46176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 45926 54622 46128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45927 86372 46128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 45876 86372 46176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 45676 86372 46376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 43876 1014 44576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 44076 27272 44376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 44126 54622 44328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 44127 86372 44328 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 44076 86372 44376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 43876 86372 44576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42076 1014 42776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42276 27272 42576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42327 86372 42528 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 42276 86372 42576 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 42076 86372 42776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40276 1014 40976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40476 27272 40776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40527 86372 40728 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 40476 86372 40776 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38727 86372 38928 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 38676 86372 38976 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36927 86372 37128 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 36876 86372 37176 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 60460 35158 86372 35298 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58791 34536 86372 35016 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 34536 86372 35326 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83360 35126 86372 35326 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 66497 26434 67739 28412 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 77297 26434 78539 28412 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28412 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 26435 86372 28416 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21826 57681 23199 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 22291 57681 23199 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61807 14328 86372 17730 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 42261 10740 86372 11491 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 10173 84482 11493 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61805 10175 84482 11491 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 6984 57736 8930 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 6984 62747 7596 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 6980 84787 7595 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61802 6981 84787 7595 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 2502 1014 3772 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 60886 3420 86372 3772 6 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 6 VSS
port 30 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 96976
string LEFclass BLOCK
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2941440
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2876172
<< end >>
