* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.inc "/import/yukari1/lrburle/OSU_180/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/OSU_180/char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL VSS

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp12t3v3__dffn_1 D Q QN CLK
X0 a_75_109 a_52_14 a_19_14 VDD pmos_3p3 w=34 l=6
X1 a_19_14 a_52_81 a_42_109 VDD pmos_3p3 w=34 l=6
X2 a_131_19 a_52_14 a_114_19 VSS nmos_3p3 w=17 l=6
X3 a_42_109 D VDD VDD pmos_3p3 w=34 l=6
X4 VDD a_19_14 a_9_19 VDD pmos_3p3 w=34 l=6
X5 a_75_19 a_52_81 a_19_14 VSS nmos_3p3 w=17 l=6
X6 VDD a_135_68 QN VDD pmos_3p3 w=34 l=6
X7 Q QN VDD VDD pmos_3p3 w=34 l=6
X8 Q QN VSS VSS nmos_3p3 w=17 l=6
X9 VSS a_135_68 a_131_19 VSS nmos_3p3 w=17 l=6
X10 a_19_14 a_52_14 a_42_19 VSS nmos_3p3 w=17 l=6
X11 VSS a_19_14 a_9_19 VSS nmos_3p3 w=17 l=6
X12 VSS a_135_68 QN VSS nmos_3p3 w=17 l=6
X13 a_52_14 a_52_81 VDD VDD pmos_3p3 w=34 l=6
X14 VDD a_135_68 a_131_109 VDD pmos_3p3 w=34 l=6
X15 VSS CLK a_52_81 VSS nmos_3p3 w=17 l=6
X16 a_131_109 a_52_81 a_114_19 VDD pmos_3p3 w=34 l=6
X17 a_114_19 a_52_14 a_103_109 VDD pmos_3p3 w=34 l=6
X18 a_135_68 a_114_19 VDD VDD pmos_3p3 w=34 l=6
X19 a_114_19 a_52_81 a_103_19 VSS nmos_3p3 w=17 l=6
X20 a_52_14 a_52_81 VSS VSS nmos_3p3 w=17 l=6
X21 a_103_109 a_9_19 VDD VDD pmos_3p3 w=34 l=6
X22 a_42_19 D VSS VSS nmos_3p3 w=17 l=6
X23 VDD a_9_19 a_75_109 VDD pmos_3p3 w=34 l=6
X24 a_103_19 a_9_19 VSS VSS nmos_3p3 w=17 l=6
X25 a_135_68 a_114_19 VSS VSS nmos_3p3 w=17 l=6
X26 VDD CLK a_52_81 VDD pmos_3p3 w=34 l=6
X27 VSS a_9_19 a_75_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
