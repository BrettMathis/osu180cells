magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 120
<< mvndiff >>
rect -88 83 0 120
rect -88 37 -75 83
rect -29 37 0 83
rect -88 0 0 37
rect 120 83 208 120
rect 120 37 149 83
rect 195 37 208 83
rect 120 0 208 37
<< mvndiffc >>
rect -75 37 -29 83
rect 149 37 195 83
<< polysilicon >>
rect 0 120 120 164
rect 0 -44 120 0
<< metal1 >>
rect -75 83 -29 120
rect -75 0 -29 37
rect 149 83 195 120
rect 149 0 195 37
<< labels >>
flabel metal1 s -52 60 -52 60 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 60 172 60 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 208112
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 207088
<< end >>
