magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect -64 1045 55 1046
rect -64 1005 64 1045
rect -64 953 -26 1005
rect 26 953 64 1005
rect -64 788 64 953
rect -64 736 -26 788
rect 26 736 64 788
rect -64 570 64 736
rect -64 518 -26 570
rect 26 518 64 570
rect -64 353 64 518
rect -64 301 -26 353
rect 26 301 64 353
rect -64 135 64 301
rect -64 83 -26 135
rect 26 83 64 135
rect -64 -83 64 83
rect -64 -135 -26 -83
rect 26 -135 64 -83
rect -64 -301 64 -135
rect -64 -353 -26 -301
rect 26 -353 64 -301
rect -64 -518 64 -353
rect -64 -570 -26 -518
rect 26 -570 64 -518
rect -64 -736 64 -570
rect -64 -788 -26 -736
rect 26 -788 64 -736
rect -64 -953 64 -788
rect -64 -1005 -26 -953
rect 26 -1005 64 -953
rect -64 -1046 64 -1005
<< via1 >>
rect -26 953 26 1005
rect -26 736 26 788
rect -26 518 26 570
rect -26 301 26 353
rect -26 83 26 135
rect -26 -135 26 -83
rect -26 -353 26 -301
rect -26 -570 26 -518
rect -26 -788 26 -736
rect -26 -1005 26 -953
<< metal2 >>
rect -64 1005 64 1045
rect -64 953 -26 1005
rect 26 953 64 1005
rect -64 788 64 953
rect -64 736 -26 788
rect 26 736 64 788
rect -64 570 64 736
rect -64 518 -26 570
rect 26 518 64 570
rect -64 353 64 518
rect -64 301 -26 353
rect 26 301 64 353
rect -64 135 64 301
rect -64 83 -26 135
rect 26 83 64 135
rect -64 -83 64 83
rect -64 -135 -26 -83
rect 26 -135 64 -83
rect -64 -301 64 -135
rect -64 -353 -26 -301
rect 26 -353 64 -301
rect -64 -518 64 -353
rect -64 -570 -26 -518
rect 26 -570 64 -518
rect -64 -736 64 -570
rect -64 -788 -26 -736
rect 26 -788 64 -736
rect -64 -953 64 -788
rect -64 -1005 -26 -953
rect 26 -1005 64 -953
rect -64 -1046 64 -1005
<< properties >>
string GDS_END 292274
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 291486
<< end >>
