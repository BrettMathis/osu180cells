* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.inc "/import/yukari1/lrburle/OSU_180/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/OSU_180/char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL VSS

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp12t3v3__dffs_1 D SN Q QN CLK
X0 a_75_109 D VDD VDD pmos_3p3 w=34 l=6
X1 Q QN VSS VSS nmos_3p3 w=17 l=6
X2 a_227_19 a_147_19 VSS VSS nmos_3p3 w=17 l=6
X3 a_208_109 SN VDD VDD pmos_3p3 w=34 l=6
X4 VSS SN a_108_19 VSS nmos_3p3 w=17 l=6
X5 VDD a_147_19 a_208_109 VDD pmos_3p3 w=34 l=6
X6 a_85_14 CLK VSS VSS nmos_3p3 w=17 l=6
X7 a_168_68 SN a_227_19 VSS nmos_3p3 w=17 l=6
X8 a_75_19 D VSS VSS nmos_3p3 w=17 l=6
X9 a_85_14 CLK VDD VDD pmos_3p3 w=34 l=6
X10 VDD a_168_68 a_164_109 VDD pmos_3p3 w=34 l=6
X11 VDD SN SN VDD pmos_3p3 w=34 l=6
X12 SN a_34_14 VDD VDD pmos_3p3 w=34 l=6
X13 a_147_19 a_85_14 a_136_109 VDD pmos_3p3 w=34 l=6
X14 a_164_109 CLK a_147_19 VDD pmos_3p3 w=34 l=6
X15 a_136_109 SN VDD VDD pmos_3p3 w=34 l=6
X16 a_136_19 SN VSS VSS nmos_3p3 w=17 l=6
X17 VDD SN a_108_109 VDD pmos_3p3 w=34 l=6
X18 VSS a_168_68 QN VSS nmos_3p3 w=17 l=6
X19 a_108_109 a_85_14 a_34_14 VDD pmos_3p3 w=34 l=6
X20 a_164_19 a_85_14 a_147_19 VSS nmos_3p3 w=17 l=6
X21 Q QN VDD VDD pmos_3p3 w=34 l=6
X22 VDD a_168_68 QN VDD pmos_3p3 w=34 l=6
X23 a_147_19 CLK a_136_19 VSS nmos_3p3 w=17 l=6
X24 VSS a_168_68 a_164_19 VSS nmos_3p3 w=17 l=6
X25 a_34_14 CLK a_75_109 VDD pmos_3p3 w=34 l=6
X26 a_29_19 SN SN VSS nmos_3p3 w=17 l=6
X27 a_34_14 a_85_14 a_75_19 VSS nmos_3p3 w=17 l=6
X28 VSS a_34_14 a_29_19 VSS nmos_3p3 w=17 l=6
X29 a_108_19 CLK a_34_14 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
