magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 2016 844
rect 297 657 365 724
rect 1313 635 1537 724
rect 1469 506 1537 635
rect 1684 468 1772 678
rect 1887 514 1955 724
rect 1684 421 1876 468
rect 186 240 671 320
rect 1786 243 1876 421
rect 1674 192 1876 243
rect 317 60 385 127
rect 1344 60 1390 138
rect 1674 106 1720 192
rect 1887 60 1955 127
rect 0 -60 2016 60
<< obsm1 >>
rect 49 481 117 621
rect 49 413 653 481
rect 49 180 95 413
rect 744 382 790 632
rect 908 493 954 632
rect 908 447 1231 493
rect 744 336 1097 382
rect 1167 371 1231 447
rect 49 134 117 180
rect 744 154 821 336
rect 1167 325 1708 371
rect 1167 211 1231 325
rect 908 143 1231 211
<< labels >>
rlabel metal1 s 186 240 671 320 6 I
port 1 nsew default input
rlabel metal1 s 1684 468 1772 678 6 Z
port 2 nsew default output
rlabel metal1 s 1684 421 1876 468 6 Z
port 2 nsew default output
rlabel metal1 s 1786 243 1876 421 6 Z
port 2 nsew default output
rlabel metal1 s 1674 192 1876 243 6 Z
port 2 nsew default output
rlabel metal1 s 1674 106 1720 192 6 Z
port 2 nsew default output
rlabel metal1 s 0 724 2016 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1887 657 1955 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1313 657 1537 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1887 635 1955 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1313 635 1537 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1887 514 1955 635 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1469 514 1537 635 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1469 506 1537 514 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1344 127 1390 138 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1887 60 1955 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1344 60 1390 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2016 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2016 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1078032
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1073628
<< end >>
