VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ffra
  CLASS BLOCK ;
  FOREIGN ffra ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 38.640 900.000 39.200 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 113.120 900.000 113.680 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 187.600 900.000 188.160 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 262.080 900.000 262.640 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 336.560 900.000 337.120 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 411.040 900.000 411.600 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 485.520 900.000 486.080 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 560.000 900.000 560.560 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 38.640 4.000 39.200 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 113.120 4.000 113.680 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 187.600 4.000 188.160 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 262.080 4.000 262.640 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 336.560 4.000 337.120 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 411.040 4.000 411.600 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 485.520 4.000 486.080 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 560.000 4.000 560.560 ;
    END
  END b[7]
  PIN ci[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 125.440 0.000 126.000 4.000 ;
    END
  END ci[0]
  PIN ci[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 623.840 0.000 624.400 4.000 ;
    END
  END ci[10]
  PIN ci[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 673.680 0.000 674.240 4.000 ;
    END
  END ci[11]
  PIN ci[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 723.520 0.000 724.080 4.000 ;
    END
  END ci[12]
  PIN ci[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 773.360 0.000 773.920 4.000 ;
    END
  END ci[13]
  PIN ci[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 823.200 0.000 823.760 4.000 ;
    END
  END ci[14]
  PIN ci[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 873.040 0.000 873.600 4.000 ;
    END
  END ci[15]
  PIN ci[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 175.280 0.000 175.840 4.000 ;
    END
  END ci[1]
  PIN ci[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END ci[2]
  PIN ci[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 274.960 0.000 275.520 4.000 ;
    END
  END ci[3]
  PIN ci[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 324.800 0.000 325.360 4.000 ;
    END
  END ci[4]
  PIN ci[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 374.640 0.000 375.200 4.000 ;
    END
  END ci[5]
  PIN ci[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 424.480 0.000 425.040 4.000 ;
    END
  END ci[6]
  PIN ci[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 474.320 0.000 474.880 4.000 ;
    END
  END ci[7]
  PIN ci[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 524.160 0.000 524.720 4.000 ;
    END
  END ci[8]
  PIN ci[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 574.000 0.000 574.560 4.000 ;
    END
  END ci[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END clk
  PIN o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 29.680 596.000 30.240 600.000 ;
    END
  END o[0]
  PIN o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 589.680 596.000 590.240 600.000 ;
    END
  END o[10]
  PIN o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 645.680 596.000 646.240 600.000 ;
    END
  END o[11]
  PIN o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 701.680 596.000 702.240 600.000 ;
    END
  END o[12]
  PIN o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 757.680 596.000 758.240 600.000 ;
    END
  END o[13]
  PIN o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 813.680 596.000 814.240 600.000 ;
    END
  END o[14]
  PIN o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 869.680 596.000 870.240 600.000 ;
    END
  END o[15]
  PIN o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 85.680 596.000 86.240 600.000 ;
    END
  END o[1]
  PIN o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 141.680 596.000 142.240 600.000 ;
    END
  END o[2]
  PIN o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 197.680 596.000 198.240 600.000 ;
    END
  END o[3]
  PIN o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 253.680 596.000 254.240 600.000 ;
    END
  END o[4]
  PIN o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 309.680 596.000 310.240 600.000 ;
    END
  END o[5]
  PIN o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 365.680 596.000 366.240 600.000 ;
    END
  END o[6]
  PIN o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 421.680 596.000 422.240 600.000 ;
    END
  END o[7]
  PIN o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 477.680 596.000 478.240 600.000 ;
    END
  END o[8]
  PIN o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 533.680 596.000 534.240 600.000 ;
    END
  END o[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 75.600 0.000 76.160 4.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET4 ;
        RECT 16.720 24.300 18.320 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 170.320 24.300 171.920 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 323.920 24.300 325.520 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 477.520 24.300 479.120 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 631.120 24.300 632.720 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 784.720 24.300 786.320 572.250 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET4 ;
        RECT 93.520 24.300 95.120 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 247.120 24.300 248.720 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 400.720 24.300 402.320 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 554.320 24.300 555.920 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 707.920 24.300 709.520 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 861.520 24.300 863.120 572.250 ;
    END
  END vss
  OBS
      LAYER MET1 ;
        RECT 1.200 24.300 898.800 572.250 ;
      LAYER MET2 ;
        RECT 3.080 595.700 29.380 596.820 ;
        RECT 30.540 595.700 85.380 596.820 ;
        RECT 86.540 595.700 141.380 596.820 ;
        RECT 142.540 595.700 197.380 596.820 ;
        RECT 198.540 595.700 253.380 596.820 ;
        RECT 254.540 595.700 309.380 596.820 ;
        RECT 310.540 595.700 365.380 596.820 ;
        RECT 366.540 595.700 421.380 596.820 ;
        RECT 422.540 595.700 477.380 596.820 ;
        RECT 478.540 595.700 533.380 596.820 ;
        RECT 534.540 595.700 589.380 596.820 ;
        RECT 590.540 595.700 645.380 596.820 ;
        RECT 646.540 595.700 701.380 596.820 ;
        RECT 702.540 595.700 757.380 596.820 ;
        RECT 758.540 595.700 813.380 596.820 ;
        RECT 814.540 595.700 869.380 596.820 ;
        RECT 870.540 595.700 898.660 596.820 ;
        RECT 3.080 4.300 898.660 595.700 ;
        RECT 3.080 4.000 25.460 4.300 ;
        RECT 26.620 4.000 75.300 4.300 ;
        RECT 76.460 4.000 125.140 4.300 ;
        RECT 126.300 4.000 174.980 4.300 ;
        RECT 176.140 4.000 224.820 4.300 ;
        RECT 225.980 4.000 274.660 4.300 ;
        RECT 275.820 4.000 324.500 4.300 ;
        RECT 325.660 4.000 374.340 4.300 ;
        RECT 375.500 4.000 424.180 4.300 ;
        RECT 425.340 4.000 474.020 4.300 ;
        RECT 475.180 4.000 523.860 4.300 ;
        RECT 525.020 4.000 573.700 4.300 ;
        RECT 574.860 4.000 623.540 4.300 ;
        RECT 624.700 4.000 673.380 4.300 ;
        RECT 674.540 4.000 723.220 4.300 ;
        RECT 724.380 4.000 773.060 4.300 ;
        RECT 774.220 4.000 822.900 4.300 ;
        RECT 824.060 4.000 872.740 4.300 ;
        RECT 873.900 4.000 898.660 4.300 ;
      LAYER MET3 ;
        RECT 4.000 560.860 898.710 572.090 ;
        RECT 4.300 559.700 895.700 560.860 ;
        RECT 4.000 486.380 898.710 559.700 ;
        RECT 4.300 485.220 895.700 486.380 ;
        RECT 4.000 411.900 898.710 485.220 ;
        RECT 4.300 410.740 895.700 411.900 ;
        RECT 4.000 337.420 898.710 410.740 ;
        RECT 4.300 336.260 895.700 337.420 ;
        RECT 4.000 262.940 898.710 336.260 ;
        RECT 4.300 261.780 895.700 262.940 ;
        RECT 4.000 188.460 898.710 261.780 ;
        RECT 4.300 187.300 895.700 188.460 ;
        RECT 4.000 113.980 898.710 187.300 ;
        RECT 4.300 112.820 895.700 113.980 ;
        RECT 4.000 39.500 898.710 112.820 ;
        RECT 4.300 38.340 895.700 39.500 ;
        RECT 4.000 24.460 898.710 38.340 ;
      LAYER MET4 ;
        RECT 32.060 263.850 93.220 378.470 ;
        RECT 95.420 263.850 170.020 378.470 ;
        RECT 172.220 263.850 246.820 378.470 ;
        RECT 249.020 263.850 323.620 378.470 ;
        RECT 325.820 263.850 400.420 378.470 ;
        RECT 402.620 263.850 477.220 378.470 ;
        RECT 479.420 263.850 554.020 378.470 ;
        RECT 556.220 263.850 630.820 378.470 ;
        RECT 633.020 263.850 706.580 378.470 ;
  END
END ffra
END LIBRARY

