magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -231 7199 78 12460
rect 4454 10445 4923 12026
<< pmos >>
rect 4516 11282 4636 11964
rect 4741 11282 4861 11964
rect 4516 10507 4636 11189
rect 4741 10507 4861 11189
<< ndiff >>
rect 656 7988 740 8007
rect 656 7754 675 7988
rect 721 7754 740 7988
rect 656 7735 740 7754
rect 1895 7988 1979 8007
rect 1895 7754 1914 7988
rect 1960 7754 1979 7988
rect 1895 7735 1979 7754
rect 3133 7988 3217 8007
rect 3133 7754 3152 7988
rect 3198 7754 3217 7988
rect 3133 7735 3217 7754
rect 4372 7988 4456 8007
rect 4372 7754 4391 7988
rect 4437 7754 4456 7988
rect 4372 7735 4456 7754
<< ndiffc >>
rect 675 7754 721 7988
rect 1914 7754 1960 7988
rect 3152 7754 3198 7988
rect 4391 7754 4437 7988
<< psubdiff >>
rect 618 5351 778 5411
rect 618 5305 675 5351
rect 721 5305 778 5351
rect 618 5245 778 5305
rect 1857 5351 2017 5411
rect 1857 5305 1914 5351
rect 1960 5305 2017 5351
rect 1857 5245 2017 5305
rect 3095 5351 3255 5411
rect 3095 5305 3152 5351
rect 3198 5305 3255 5351
rect 3095 5245 3255 5305
rect -51 583 33 602
rect -51 443 -32 583
rect 14 443 33 583
rect -51 424 33 443
rect 1276 583 1360 602
rect 1276 443 1295 583
rect 1341 443 1360 583
rect 1276 424 1360 443
rect 2515 583 2599 602
rect 2515 443 2534 583
rect 2580 443 2599 583
rect 2515 424 2599 443
rect 3753 583 3837 602
rect 3753 443 3772 583
rect 3818 443 3837 583
rect 3753 424 3837 443
rect 4992 583 5076 602
rect 4992 443 5011 583
rect 5057 443 5076 583
rect 4992 424 5076 443
<< psubdiffcont >>
rect 675 5305 721 5351
rect 1914 5305 1960 5351
rect 3152 5305 3198 5351
rect -32 443 14 583
rect 1295 443 1341 583
rect 2534 443 2580 583
rect 3772 443 3818 583
rect 5011 443 5057 583
<< metal1 >>
rect -23 10362 4966 10436
rect 660 8015 736 8027
rect 660 7755 672 8015
rect 724 7755 736 8015
rect 660 7754 675 7755
rect 721 7754 736 7755
rect 660 7743 736 7754
rect 1899 8015 1975 8027
rect 1899 7755 1911 8015
rect 1963 7755 1975 8015
rect 1899 7754 1914 7755
rect 1960 7754 1975 7755
rect 1899 7743 1975 7754
rect 3137 8015 3213 8027
rect 3137 7755 3149 8015
rect 3201 7755 3213 8015
rect 3137 7754 3152 7755
rect 3198 7754 3213 7755
rect 3137 7743 3213 7754
rect 4376 8015 4452 8027
rect 4376 7755 4388 8015
rect 4440 7755 4452 8015
rect 4376 7754 4391 7755
rect 4437 7754 4452 7755
rect 4376 7743 4452 7754
rect 627 5351 769 5402
rect 627 5305 675 5351
rect 721 5305 769 5351
rect 627 5254 769 5305
rect 1866 5351 2008 5402
rect 1866 5305 1914 5351
rect 1960 5305 2008 5351
rect 1866 5254 2008 5305
rect 3104 5351 3246 5402
rect 3104 5305 3152 5351
rect 3198 5305 3246 5351
rect 3104 5254 3246 5305
rect 1134 1509 1210 1521
rect 1134 1457 1146 1509
rect 1198 1457 1210 1509
rect 1134 1445 1210 1457
rect 1425 1509 1501 1521
rect 1425 1457 1437 1509
rect 1489 1457 1501 1509
rect 1425 1445 1501 1457
rect 2373 1509 2449 1521
rect 2373 1457 2385 1509
rect 2437 1457 2449 1509
rect 2373 1445 2449 1457
rect 2664 1509 2740 1521
rect 2664 1457 2676 1509
rect 2728 1457 2740 1509
rect 2664 1445 2740 1457
rect 3611 1509 3687 1521
rect 3611 1457 3623 1509
rect 3675 1457 3687 1509
rect 3611 1445 3687 1457
rect 3902 1509 3978 1521
rect 3902 1457 3914 1509
rect 3966 1457 3978 1509
rect 3902 1445 3978 1457
rect -43 591 25 594
rect -43 583 68 591
rect -43 443 -32 583
rect 14 443 68 583
rect -43 90 68 443
rect 1284 583 1352 594
rect 1284 443 1295 583
rect 1341 443 1352 583
rect 1284 432 1352 443
rect 2523 583 2591 594
rect 2523 443 2534 583
rect 2580 443 2591 583
rect 2523 432 2591 443
rect 3761 583 3829 594
rect 3761 443 3772 583
rect 3818 443 3829 583
rect 3761 432 3829 443
rect 5000 583 5068 594
rect 5000 443 5011 583
rect 5057 443 5068 583
rect 5000 432 5068 443
<< via1 >>
rect 672 7988 724 8015
rect 672 7755 675 7988
rect 675 7755 721 7988
rect 721 7755 724 7988
rect 1911 7988 1963 8015
rect 1911 7755 1914 7988
rect 1914 7755 1960 7988
rect 1960 7755 1963 7988
rect 3149 7988 3201 8015
rect 3149 7755 3152 7988
rect 3152 7755 3198 7988
rect 3198 7755 3201 7988
rect 4388 7988 4440 8015
rect 4388 7755 4391 7988
rect 4391 7755 4437 7988
rect 4437 7755 4440 7988
rect 1146 1457 1198 1509
rect 1437 1457 1489 1509
rect 2385 1457 2437 1509
rect 2676 1457 2728 1509
rect 3623 1457 3675 1509
rect 3914 1457 3966 1509
<< metal2 >>
rect 660 8017 736 8027
rect 660 7753 670 8017
rect 726 7753 736 8017
rect 660 7743 736 7753
rect 1899 8017 1975 8027
rect 1899 7753 1909 8017
rect 1965 7753 1975 8017
rect 1899 7743 1975 7753
rect 3137 8017 3213 8027
rect 3137 7753 3147 8017
rect 3203 7753 3213 8017
rect 3137 7743 3213 7753
rect 4376 8017 4452 8027
rect 4376 7753 4386 8017
rect 4442 7753 4452 8017
rect 4376 7743 4452 7753
rect 1134 1511 1210 1533
rect 1134 1351 1144 1511
rect 1200 1351 1210 1511
rect 1134 1251 1210 1351
rect 1425 1511 1501 1533
rect 1425 1351 1435 1511
rect 1491 1351 1501 1511
rect 1425 1251 1501 1351
rect 2373 1511 2449 1533
rect 2373 1351 2383 1511
rect 2439 1351 2449 1511
rect 2373 1251 2449 1351
rect 2664 1511 2740 1533
rect 2664 1351 2674 1511
rect 2730 1351 2740 1511
rect 2664 1251 2740 1351
rect 3611 1511 3687 1533
rect 3611 1351 3621 1511
rect 3677 1351 3687 1511
rect 3611 1251 3687 1351
rect 3902 1511 3978 1533
rect 3902 1351 3912 1511
rect 3968 1351 3978 1511
rect 3902 1251 3978 1351
<< via2 >>
rect 670 8015 726 8017
rect 670 7755 672 8015
rect 672 7755 724 8015
rect 724 7755 726 8015
rect 670 7753 726 7755
rect 1909 8015 1965 8017
rect 1909 7755 1911 8015
rect 1911 7755 1963 8015
rect 1963 7755 1965 8015
rect 1909 7753 1965 7755
rect 3147 8015 3203 8017
rect 3147 7755 3149 8015
rect 3149 7755 3201 8015
rect 3201 7755 3203 8015
rect 3147 7753 3203 7755
rect 4386 8015 4442 8017
rect 4386 7755 4388 8015
rect 4388 7755 4440 8015
rect 4440 7755 4442 8015
rect 4386 7753 4442 7755
rect 1144 1509 1200 1511
rect 1144 1457 1146 1509
rect 1146 1457 1198 1509
rect 1198 1457 1200 1509
rect 1144 1351 1200 1457
rect 1435 1509 1491 1511
rect 1435 1457 1437 1509
rect 1437 1457 1489 1509
rect 1489 1457 1491 1509
rect 1435 1351 1491 1457
rect 2383 1509 2439 1511
rect 2383 1457 2385 1509
rect 2385 1457 2437 1509
rect 2437 1457 2439 1509
rect 2383 1351 2439 1457
rect 2674 1509 2730 1511
rect 2674 1457 2676 1509
rect 2676 1457 2728 1509
rect 2728 1457 2730 1509
rect 2674 1351 2730 1457
rect 3621 1509 3677 1511
rect 3621 1457 3623 1509
rect 3623 1457 3675 1509
rect 3675 1457 3677 1509
rect 3621 1351 3677 1457
rect 3912 1509 3968 1511
rect 3912 1457 3914 1509
rect 3914 1457 3966 1509
rect 3966 1457 3968 1509
rect 3912 1351 3968 1457
<< metal3 >>
rect -822 8017 7080 8027
rect -822 7753 670 8017
rect 726 7753 1909 8017
rect 1965 7753 3147 8017
rect 3203 7753 4386 8017
rect 4442 7753 7080 8017
rect -822 7743 7080 7753
rect 1134 1511 1210 1521
rect 1134 1351 1144 1511
rect 1200 1351 1210 1511
rect 1134 1341 1210 1351
rect 1425 1511 1501 1521
rect 1425 1351 1435 1511
rect 1491 1351 1501 1511
rect 1425 1341 1501 1351
rect 2373 1511 2449 1521
rect 2373 1351 2383 1511
rect 2439 1351 2449 1511
rect 2373 1341 2449 1351
rect 2664 1511 2740 1521
rect 2664 1351 2674 1511
rect 2730 1351 2740 1511
rect 2664 1341 2740 1351
rect 3611 1511 3687 1521
rect 3611 1351 3621 1511
rect 3677 1351 3687 1511
rect 3611 1341 3687 1351
rect 3902 1511 3978 1521
rect 3902 1351 3912 1511
rect 3968 1351 3978 1511
rect 3902 1341 3978 1351
use M1_NACTIVE4310589983232_64x8m81  M1_NACTIVE4310589983232_64x8m81_0
timestamp 1669390400
transform 1 0 1937 0 1 7871
box 0 0 1 1
use M1_NACTIVE4310589983232_64x8m81  M1_NACTIVE4310589983232_64x8m81_1
timestamp 1669390400
transform 1 0 4414 0 1 7871
box 0 0 1 1
use M1_NACTIVE4310589983232_64x8m81  M1_NACTIVE4310589983232_64x8m81_2
timestamp 1669390400
transform 1 0 3175 0 1 7871
box 0 0 1 1
use M1_NACTIVE4310589983232_64x8m81  M1_NACTIVE4310589983232_64x8m81_3
timestamp 1669390400
transform 1 0 698 0 1 7871
box 0 0 1 1
use M1_PACTIVE4310589983231_64x8m81  M1_PACTIVE4310589983231_64x8m81_0
timestamp 1669390400
transform 1 0 1318 0 1 513
box 0 0 1 1
use M1_PACTIVE4310589983231_64x8m81  M1_PACTIVE4310589983231_64x8m81_1
timestamp 1669390400
transform 1 0 2557 0 1 513
box 0 0 1 1
use M1_PACTIVE4310589983231_64x8m81  M1_PACTIVE4310589983231_64x8m81_2
timestamp 1669390400
transform 1 0 5034 0 1 513
box 0 0 1 1
use M1_PACTIVE4310589983231_64x8m81  M1_PACTIVE4310589983231_64x8m81_3
timestamp 1669390400
transform 1 0 3795 0 1 513
box 0 0 1 1
use M1_PACTIVE4310589983231_64x8m81  M1_PACTIVE4310589983231_64x8m81_4
timestamp 1669390400
transform 1 0 -9 0 1 513
box 0 0 1 1
use M1_PSUB$$45111340_64x8m81  M1_PSUB$$45111340_64x8m81_0
timestamp 1669390400
transform 1 0 1937 0 1 5328
box 0 0 1 1
use M1_PSUB$$45111340_64x8m81  M1_PSUB$$45111340_64x8m81_1
timestamp 1669390400
transform 1 0 698 0 1 5328
box 0 0 1 1
use M1_PSUB$$45111340_64x8m81  M1_PSUB$$45111340_64x8m81_2
timestamp 1669390400
transform 1 0 3175 0 1 5328
box 0 0 1 1
use M2_M14310589983228_64x8m81  M2_M14310589983228_64x8m81_0
timestamp 1669390400
transform 1 0 1463 0 1 1483
box 0 0 1 1
use M2_M14310589983228_64x8m81  M2_M14310589983228_64x8m81_1
timestamp 1669390400
transform 1 0 2702 0 1 1483
box 0 0 1 1
use M2_M14310589983228_64x8m81  M2_M14310589983228_64x8m81_2
timestamp 1669390400
transform 1 0 2411 0 1 1483
box 0 0 1 1
use M2_M14310589983228_64x8m81  M2_M14310589983228_64x8m81_3
timestamp 1669390400
transform 1 0 3940 0 1 1483
box 0 0 1 1
use M2_M14310589983228_64x8m81  M2_M14310589983228_64x8m81_4
timestamp 1669390400
transform 1 0 3649 0 1 1483
box 0 0 1 1
use M2_M14310589983228_64x8m81  M2_M14310589983228_64x8m81_5
timestamp 1669390400
transform 1 0 1172 0 1 1483
box 0 0 1 1
use M2_M14310589983233_64x8m81  M2_M14310589983233_64x8m81_0
timestamp 1669390400
transform 1 0 1937 0 1 7885
box 0 0 1 1
use M2_M14310589983233_64x8m81  M2_M14310589983233_64x8m81_1
timestamp 1669390400
transform 1 0 3175 0 1 7885
box 0 0 1 1
use M2_M14310589983233_64x8m81  M2_M14310589983233_64x8m81_2
timestamp 1669390400
transform 1 0 4414 0 1 7885
box 0 0 1 1
use M2_M14310589983233_64x8m81  M2_M14310589983233_64x8m81_3
timestamp 1669390400
transform 1 0 698 0 1 7885
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_0
timestamp 1669390400
transform 1 0 1463 0 1 1431
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_1
timestamp 1669390400
transform 1 0 2411 0 1 1431
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_2
timestamp 1669390400
transform 1 0 2702 0 1 1431
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_3
timestamp 1669390400
transform 1 0 3649 0 1 1431
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_4
timestamp 1669390400
transform 1 0 3940 0 1 1431
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_5
timestamp 1669390400
transform 1 0 1172 0 1 1431
box 0 0 1 1
use M3_M24310589983230_64x8m81  M3_M24310589983230_64x8m81_0
timestamp 1669390400
transform 1 0 698 0 1 7885
box 0 0 1 1
use M3_M24310589983230_64x8m81  M3_M24310589983230_64x8m81_1
timestamp 1669390400
transform 1 0 3175 0 1 7885
box 0 0 1 1
use M3_M24310589983230_64x8m81  M3_M24310589983230_64x8m81_2
timestamp 1669390400
transform 1 0 4414 0 1 7885
box 0 0 1 1
use M3_M24310589983230_64x8m81  M3_M24310589983230_64x8m81_3
timestamp 1669390400
transform 1 0 1937 0 1 7885
box 0 0 1 1
use ypass_gate_64x8m81  ypass_gate_64x8m81_0
timestamp 1669390400
transform -1 0 3175 0 1 91
box -221 -10 930 12370
use ypass_gate_64x8m81  ypass_gate_64x8m81_1
timestamp 1669390400
transform -1 0 4414 0 1 91
box -221 -10 930 12370
use ypass_gate_64x8m81  ypass_gate_64x8m81_2
timestamp 1669390400
transform -1 0 1937 0 1 91
box -221 -10 930 12370
use ypass_gate_64x8m81  ypass_gate_64x8m81_3
timestamp 1669390400
transform -1 0 698 0 1 91
box -221 -10 930 12370
use ypass_gate_64x8m81  ypass_gate_64x8m81_4
timestamp 1669390400
transform 1 0 3175 0 1 91
box -221 -10 930 12370
use ypass_gate_64x8m81  ypass_gate_64x8m81_5
timestamp 1669390400
transform 1 0 1937 0 1 91
box -221 -10 930 12370
use ypass_gate_64x8m81  ypass_gate_64x8m81_6
timestamp 1669390400
transform 1 0 698 0 1 91
box -221 -10 930 12370
use ypass_gate_a_64x8m81  ypass_gate_a_64x8m81_0
timestamp 1669390400
transform 1 0 4414 0 1 91
box -221 -10 787 12370
<< properties >>
string GDS_END 581262
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 577850
<< end >>
