magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 408 300
<< mvpmos >>
rect 0 0 200 180
<< mvpdiff >>
rect -88 167 0 180
rect -88 121 -75 167
rect -29 121 0 167
rect -88 59 0 121
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 200 167 288 180
rect 200 121 229 167
rect 275 121 288 167
rect 200 59 288 121
rect 200 13 229 59
rect 275 13 288 59
rect 200 0 288 13
<< mvpdiffc >>
rect -75 121 -29 167
rect -75 13 -29 59
rect 229 121 275 167
rect 229 13 275 59
<< polysilicon >>
rect 0 180 200 224
rect 0 -44 200 0
<< metal1 >>
rect -75 167 -29 180
rect -75 59 -29 121
rect -75 0 -29 13
rect 229 167 275 180
rect 229 59 275 121
rect 229 0 275 13
<< labels >>
flabel metal1 s -52 90 -52 90 0 FreeSans 400 0 0 0 S
flabel metal1 s 252 90 252 90 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 637068
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 635852
<< end >>
