magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 3558 1094
<< pwell >>
rect -86 -86 3558 453
<< mvnmos >>
rect 162 175 282 333
rect 386 175 506 333
rect 754 168 874 286
rect 1044 168 1164 286
rect 1268 168 1388 286
rect 1436 168 1556 286
rect 1660 168 1780 286
rect 1928 215 2048 333
rect 2152 215 2272 333
rect 2412 69 2532 333
rect 2636 69 2756 333
rect 3004 69 3124 333
rect 3228 69 3348 333
<< mvpmos >>
rect 202 573 302 849
rect 406 573 506 849
rect 774 593 874 793
rect 978 593 1078 793
rect 1268 593 1368 793
rect 1456 593 1556 793
rect 1660 593 1760 793
rect 1864 593 1964 793
rect 2180 593 2280 793
rect 2432 573 2532 939
rect 2636 573 2736 939
rect 3035 573 3135 939
rect 3239 573 3339 939
<< mvndiff >>
rect 74 320 162 333
rect 74 274 87 320
rect 133 274 162 320
rect 74 175 162 274
rect 282 234 386 333
rect 282 188 311 234
rect 357 188 386 234
rect 282 175 386 188
rect 506 320 594 333
rect 506 274 535 320
rect 581 274 594 320
rect 1840 320 1928 333
rect 1840 286 1853 320
rect 506 175 594 274
rect 666 227 754 286
rect 666 181 679 227
rect 725 181 754 227
rect 666 168 754 181
rect 874 273 1044 286
rect 874 227 912 273
rect 958 227 1044 273
rect 874 168 1044 227
rect 1164 273 1268 286
rect 1164 227 1193 273
rect 1239 227 1268 273
rect 1164 168 1268 227
rect 1388 168 1436 286
rect 1556 227 1660 286
rect 1556 181 1585 227
rect 1631 181 1660 227
rect 1556 168 1660 181
rect 1780 274 1853 286
rect 1899 274 1928 320
rect 1780 215 1928 274
rect 2048 320 2152 333
rect 2048 274 2077 320
rect 2123 274 2152 320
rect 2048 215 2152 274
rect 2272 320 2412 333
rect 2272 274 2337 320
rect 2383 274 2412 320
rect 2272 215 2412 274
rect 1780 168 1860 215
rect 2332 69 2412 215
rect 2532 222 2636 333
rect 2532 82 2561 222
rect 2607 82 2636 222
rect 2532 69 2636 82
rect 2756 320 2844 333
rect 2756 274 2785 320
rect 2831 274 2844 320
rect 2756 69 2844 274
rect 2916 128 3004 333
rect 2916 82 2929 128
rect 2975 82 3004 128
rect 2916 69 3004 82
rect 3124 320 3228 333
rect 3124 274 3153 320
rect 3199 274 3228 320
rect 3124 69 3228 274
rect 3348 222 3436 333
rect 3348 82 3377 222
rect 3423 82 3436 222
rect 3348 69 3436 82
<< mvpdiff >>
rect 114 739 202 849
rect 114 599 127 739
rect 173 599 202 739
rect 114 573 202 599
rect 302 836 406 849
rect 302 696 331 836
rect 377 696 406 836
rect 302 573 406 696
rect 506 632 594 849
rect 2352 793 2432 939
rect 506 586 535 632
rect 581 586 594 632
rect 686 780 774 793
rect 686 734 699 780
rect 745 734 774 780
rect 686 593 774 734
rect 874 746 978 793
rect 874 606 903 746
rect 949 606 978 746
rect 874 593 978 606
rect 1078 746 1268 793
rect 1078 606 1193 746
rect 1239 606 1268 746
rect 1078 593 1268 606
rect 1368 593 1456 793
rect 1556 780 1660 793
rect 1556 640 1585 780
rect 1631 640 1660 780
rect 1556 593 1660 640
rect 1760 746 1864 793
rect 1760 606 1789 746
rect 1835 606 1864 746
rect 1760 593 1864 606
rect 1964 746 2180 793
rect 1964 606 2077 746
rect 2123 606 2180 746
rect 1964 593 2180 606
rect 2280 773 2432 793
rect 2280 633 2357 773
rect 2403 633 2432 773
rect 2280 593 2432 633
rect 506 573 594 586
rect 2352 573 2432 593
rect 2532 926 2636 939
rect 2532 880 2561 926
rect 2607 880 2636 926
rect 2532 573 2636 880
rect 2736 632 2824 939
rect 2736 586 2765 632
rect 2811 586 2824 632
rect 2736 573 2824 586
rect 2947 926 3035 939
rect 2947 880 2960 926
rect 3006 880 3035 926
rect 2947 573 3035 880
rect 3135 632 3239 939
rect 3135 586 3164 632
rect 3210 586 3239 632
rect 3135 573 3239 586
rect 3339 926 3427 939
rect 3339 786 3368 926
rect 3414 786 3427 926
rect 3339 573 3427 786
<< mvndiffc >>
rect 87 274 133 320
rect 311 188 357 234
rect 535 274 581 320
rect 679 181 725 227
rect 912 227 958 273
rect 1193 227 1239 273
rect 1585 181 1631 227
rect 1853 274 1899 320
rect 2077 274 2123 320
rect 2337 274 2383 320
rect 2561 82 2607 222
rect 2785 274 2831 320
rect 2929 82 2975 128
rect 3153 274 3199 320
rect 3377 82 3423 222
<< mvpdiffc >>
rect 127 599 173 739
rect 331 696 377 836
rect 535 586 581 632
rect 699 734 745 780
rect 903 606 949 746
rect 1193 606 1239 746
rect 1585 640 1631 780
rect 1789 606 1835 746
rect 2077 606 2123 746
rect 2357 633 2403 773
rect 2561 880 2607 926
rect 2765 586 2811 632
rect 2960 880 3006 926
rect 3164 586 3210 632
rect 3368 786 3414 926
<< polysilicon >>
rect 406 909 1078 949
rect 2432 939 2532 983
rect 2636 939 2736 983
rect 3035 939 3135 983
rect 3239 939 3339 983
rect 202 849 302 893
rect 406 849 506 909
rect 774 793 874 837
rect 978 793 1078 909
rect 1268 885 1964 925
rect 1268 872 1368 885
rect 1268 826 1281 872
rect 1327 826 1368 872
rect 1268 793 1368 826
rect 1456 793 1556 837
rect 1660 793 1760 837
rect 1864 793 1964 885
rect 2180 793 2280 837
rect 202 523 302 573
rect 202 477 215 523
rect 261 477 302 523
rect 202 393 302 477
rect 406 412 506 573
rect 162 333 282 393
rect 406 377 419 412
rect 386 366 419 377
rect 465 366 506 412
rect 386 333 506 366
rect 774 413 874 593
rect 978 549 1078 593
rect 1268 533 1368 593
rect 774 367 814 413
rect 860 367 874 413
rect 774 330 874 367
rect 1124 493 1368 533
rect 1456 560 1556 593
rect 1456 514 1497 560
rect 1543 514 1556 560
rect 1124 330 1164 493
rect 754 286 874 330
rect 1044 286 1164 330
rect 1268 365 1388 378
rect 1268 319 1329 365
rect 1375 319 1388 365
rect 1456 330 1556 514
rect 1268 286 1388 319
rect 1436 286 1556 330
rect 1660 468 1760 593
rect 1660 422 1673 468
rect 1719 422 1760 468
rect 1864 501 1964 593
rect 2180 549 2280 593
rect 1864 461 2192 501
rect 1660 330 1760 422
rect 2152 377 2192 461
rect 2240 497 2280 549
rect 2240 484 2312 497
rect 2240 438 2253 484
rect 2299 438 2312 484
rect 2240 425 2312 438
rect 2432 430 2532 573
rect 2432 384 2473 430
rect 2519 384 2532 430
rect 2432 377 2532 384
rect 1928 333 2048 377
rect 2152 333 2272 377
rect 2412 333 2532 377
rect 2636 540 2736 573
rect 2636 494 2649 540
rect 2695 494 2736 540
rect 2636 377 2736 494
rect 3035 465 3135 573
rect 3239 465 3339 573
rect 3004 412 3339 465
rect 2636 333 2756 377
rect 3004 366 3048 412
rect 3094 393 3339 412
rect 3094 366 3124 393
rect 3004 333 3124 366
rect 3228 377 3339 393
rect 3228 333 3348 377
rect 1660 286 1780 330
rect 162 131 282 175
rect 386 76 506 175
rect 1928 182 2048 215
rect 754 124 874 168
rect 1044 124 1164 168
rect 1268 76 1388 168
rect 1436 124 1556 168
rect 1660 124 1780 168
rect 1928 136 1941 182
rect 1987 136 2048 182
rect 2152 171 2272 215
rect 1928 123 2048 136
rect 386 36 1388 76
rect 2412 25 2532 69
rect 2636 25 2756 69
rect 3004 25 3124 69
rect 3228 25 3348 69
<< polycontact >>
rect 1281 826 1327 872
rect 215 477 261 523
rect 419 366 465 412
rect 814 367 860 413
rect 1497 514 1543 560
rect 1329 319 1375 365
rect 1673 422 1719 468
rect 2253 438 2299 484
rect 2473 384 2519 430
rect 2649 494 2695 540
rect 3048 366 3094 412
rect 1941 136 1987 182
<< metal1 >>
rect 0 926 3472 1098
rect 0 918 2561 926
rect 331 836 377 918
rect 127 739 173 750
rect 699 780 745 918
rect 699 723 745 734
rect 791 826 1281 872
rect 1327 826 1338 872
rect 331 685 377 696
rect 791 643 837 826
rect 1585 780 1631 918
rect 2607 918 2960 926
rect 2561 869 2607 880
rect 3006 918 3368 926
rect 2960 869 3006 880
rect 3414 918 3472 926
rect 173 599 465 634
rect 127 588 465 599
rect 142 523 373 542
rect 142 477 215 523
rect 261 477 373 523
rect 142 466 373 477
rect 419 412 465 588
rect 419 348 465 366
rect 87 320 465 348
rect 133 302 465 320
rect 535 632 837 643
rect 581 597 837 632
rect 903 746 958 757
rect 949 606 958 746
rect 903 595 958 606
rect 535 320 581 586
rect 680 413 865 447
rect 680 367 814 413
rect 860 367 865 413
rect 680 338 865 367
rect 87 263 133 274
rect 535 263 581 274
rect 912 273 958 595
rect 311 234 357 245
rect 311 90 357 188
rect 679 227 725 238
rect 912 216 958 227
rect 1193 746 1239 757
rect 2357 773 3310 784
rect 3368 775 3414 786
rect 1585 629 1631 640
rect 1789 746 1835 757
rect 1193 457 1239 606
rect 1789 571 1835 606
rect 1497 560 1835 571
rect 1543 525 1835 560
rect 1497 503 1543 514
rect 1673 468 1719 479
rect 1193 422 1673 457
rect 1193 411 1719 422
rect 1789 457 1835 525
rect 2077 746 2123 757
rect 2403 738 3310 773
rect 2357 622 2403 633
rect 2765 632 2811 643
rect 2077 576 2123 606
rect 2077 540 2706 576
rect 2077 530 2649 540
rect 1789 411 1899 457
rect 1193 273 1239 411
rect 1318 319 1329 365
rect 1375 319 1807 365
rect 1193 216 1239 227
rect 1585 227 1631 238
rect 679 90 725 181
rect 1585 90 1631 181
rect 1761 182 1807 319
rect 1853 320 1899 411
rect 1853 263 1899 274
rect 2077 320 2123 530
rect 2638 494 2649 530
rect 2695 494 2706 540
rect 2077 263 2123 274
rect 2234 438 2253 484
rect 2299 438 2310 484
rect 2234 182 2280 438
rect 2765 430 2811 586
rect 2462 384 2473 430
rect 2519 412 2811 430
rect 3164 632 3218 654
rect 3210 586 3218 632
rect 2519 384 3048 412
rect 2774 366 3048 384
rect 3094 366 3105 412
rect 2326 320 2728 325
rect 2326 274 2337 320
rect 2383 279 2728 320
rect 2383 274 2394 279
rect 1761 136 1941 182
rect 1987 136 2280 182
rect 2561 222 2607 233
rect 0 82 2561 90
rect 2682 228 2728 279
rect 2774 320 2842 366
rect 3164 320 3218 586
rect 2774 274 2785 320
rect 2831 274 2842 320
rect 3142 274 3153 320
rect 3199 274 3218 320
rect 3264 228 3310 738
rect 2682 182 3310 228
rect 3377 222 3423 233
rect 2918 90 2929 128
rect 2607 82 2929 90
rect 2975 90 2986 128
rect 2975 82 3377 90
rect 3423 82 3472 90
rect 0 -90 3472 82
<< labels >>
flabel metal1 s 142 466 373 542 0 FreeSans 200 0 0 0 CLKN
port 2 nsew clock input
flabel metal1 s 680 338 865 447 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3164 320 3218 654 0 FreeSans 200 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 918 3472 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 311 238 357 245 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3142 274 3218 320 1 Q
port 3 nsew default output
rlabel metal1 s 3368 869 3414 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2960 869 3006 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2561 869 2607 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1585 869 1631 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 699 869 745 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 331 869 377 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3368 775 3414 869 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1585 775 1631 869 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 699 775 745 869 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 331 775 377 869 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1585 723 1631 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 699 723 745 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 331 723 377 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1585 685 1631 723 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 331 685 377 723 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1585 629 1631 685 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1585 233 1631 238 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 679 233 725 238 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 311 233 357 238 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3377 128 3423 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2561 128 2607 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1585 128 1631 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 679 128 725 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 311 128 357 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3377 90 3423 128 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2918 90 2986 128 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2561 90 2607 128 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1585 90 1631 128 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 679 90 725 128 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 311 90 357 128 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3472 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3472 1008
string GDS_END 1472818
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1464892
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
