magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< mvnmos >>
rect 0 0 120 1700
rect 224 0 344 1700
<< mvndiff >>
rect -88 1687 0 1700
rect -88 13 -75 1687
rect -29 13 0 1687
rect -88 0 0 13
rect 120 1687 224 1700
rect 120 13 149 1687
rect 195 13 224 1687
rect 120 0 224 13
rect 344 1687 432 1700
rect 344 13 373 1687
rect 419 13 432 1687
rect 344 0 432 13
<< mvndiffc >>
rect -75 13 -29 1687
rect 149 13 195 1687
rect 373 13 419 1687
<< polysilicon >>
rect 0 1700 120 1744
rect 224 1700 344 1744
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 1687 -29 1700
rect -75 0 -29 13
rect 149 1687 195 1700
rect 149 0 195 13
rect 373 1687 419 1700
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 850 -52 850 0 FreeSans 200 0 0 0 S
flabel metal1 s 396 850 396 850 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 850 172 850 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 914600
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 910058
<< end >>
