magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -208 -120 328 360
<< mvpmos >>
rect 0 0 120 240
<< mvpdiff >>
rect -88 227 0 240
rect -88 181 -75 227
rect -29 181 0 227
rect -88 59 0 181
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 227 208 240
rect 120 181 149 227
rect 195 181 208 227
rect 120 59 208 181
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvpdiffc >>
rect -75 181 -29 227
rect -75 13 -29 59
rect 149 181 195 227
rect 149 13 195 59
<< polysilicon >>
rect 0 240 120 284
rect 0 -44 120 0
<< metal1 >>
rect -75 227 -29 240
rect -75 59 -29 181
rect -75 0 -29 13
rect 149 227 195 240
rect 149 59 195 181
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 120 -52 120 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 120 172 120 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 260258
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 259042
<< end >>
