magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< polysilicon >>
rect 751 7051 871 7092
rect 1265 7051 1385 7167
rect 465 7005 871 7051
rect 465 6959 539 7005
rect 585 6959 697 7005
rect 743 6959 871 7005
rect 465 6913 871 6959
rect 975 7005 1385 7051
rect 975 6959 1049 7005
rect 1095 6959 1207 7005
rect 1253 6959 1385 7005
rect 975 6913 1385 6959
rect 751 6820 871 6913
rect 1265 5957 1385 6913
<< polycontact >>
rect 539 6959 585 7005
rect 697 6959 743 7005
rect 1049 6959 1095 7005
rect 1207 6959 1253 7005
<< metal1 >>
rect 324 8301 756 8430
rect 324 8249 459 8301
rect 511 8249 666 8301
rect 718 8249 756 8301
rect 324 8083 756 8249
rect 324 8031 459 8083
rect 511 8031 666 8083
rect 718 8031 756 8083
rect 324 7865 756 8031
rect 324 7813 459 7865
rect 511 7813 666 7865
rect 718 7813 756 7865
rect 324 7647 756 7813
rect 324 7595 459 7647
rect 511 7595 666 7647
rect 718 7595 756 7647
rect 324 7131 756 7595
rect 1148 8278 1276 8318
rect 1148 8226 1186 8278
rect 1238 8226 1276 8278
rect 1148 8060 1276 8226
rect 1148 8008 1186 8060
rect 1238 8008 1276 8060
rect 1148 7842 1276 8008
rect 1148 7790 1186 7842
rect 1238 7790 1276 7842
rect 1148 7624 1276 7790
rect 1148 7572 1186 7624
rect 1238 7572 1276 7624
rect 1148 7532 1276 7572
rect 421 7042 761 7049
rect 865 7042 980 7192
rect 421 7008 778 7042
rect 421 6956 459 7008
rect 511 7005 671 7008
rect 723 7005 778 7008
rect 511 6959 539 7005
rect 585 6959 671 7005
rect 743 6959 778 7005
rect 511 6956 671 6959
rect 723 6956 778 6959
rect 421 6922 778 6956
rect 865 7005 1288 7042
rect 865 6959 1049 7005
rect 1095 6959 1207 7005
rect 1253 6959 1288 7005
rect 865 6922 1288 6959
rect 421 6916 761 6922
rect 276 3273 756 6793
rect 865 6455 980 6922
rect 1414 5485 1460 7308
rect 1374 4490 1498 4530
rect 1374 4438 1410 4490
rect 1462 4438 1498 4490
rect 1374 4272 1498 4438
rect 1374 4220 1410 4272
rect 1462 4220 1498 4272
rect 1374 4180 1498 4220
rect 860 3583 984 3623
rect 860 3531 896 3583
rect 948 3531 984 3583
rect 860 3365 984 3531
rect 860 3313 896 3365
rect 948 3313 984 3365
rect 860 3273 984 3313
rect -106 3078 1760 3170
rect -106 2876 1760 2969
rect -106 2674 1760 2767
rect -106 2472 1760 2565
rect 423 1624 547 1664
rect 423 1572 459 1624
rect 511 1572 547 1624
rect 423 1406 547 1572
rect 423 1354 459 1406
rect 511 1354 547 1406
rect 423 1314 547 1354
<< via1 >>
rect 459 8249 511 8301
rect 666 8249 718 8301
rect 459 8031 511 8083
rect 666 8031 718 8083
rect 459 7813 511 7865
rect 666 7813 718 7865
rect 459 7595 511 7647
rect 666 7595 718 7647
rect 1186 8226 1238 8278
rect 1186 8008 1238 8060
rect 1186 7790 1238 7842
rect 1186 7572 1238 7624
rect 459 6956 511 7008
rect 671 7005 723 7008
rect 671 6959 697 7005
rect 697 6959 723 7005
rect 671 6956 723 6959
rect 1410 4438 1462 4490
rect 1410 4220 1462 4272
rect 896 3531 948 3583
rect 896 3313 948 3365
rect 459 1572 511 1624
rect 459 1354 511 1406
<< metal2 >>
rect 421 8303 756 8341
rect 421 8247 457 8303
rect 513 8247 664 8303
rect 720 8247 756 8303
rect 421 8085 756 8247
rect 421 8029 457 8085
rect 513 8029 664 8085
rect 720 8029 756 8085
rect 421 7867 756 8029
rect 421 7811 457 7867
rect 513 7811 664 7867
rect 720 7811 756 7867
rect 421 7649 756 7811
rect 421 7593 457 7649
rect 513 7593 664 7649
rect 720 7593 756 7649
rect 421 7555 756 7593
rect 1148 8280 1276 8317
rect 1148 8224 1184 8280
rect 1240 8224 1276 8280
rect 1148 8062 1276 8224
rect 1148 8006 1184 8062
rect 1240 8006 1276 8062
rect 1148 7844 1276 8006
rect 1148 7788 1184 7844
rect 1240 7788 1276 7844
rect 1148 7626 1276 7788
rect 1148 7570 1184 7626
rect 1240 7570 1276 7626
rect 1148 7532 1276 7570
rect 421 7008 761 7049
rect 421 6956 459 7008
rect 511 6956 671 7008
rect 723 6956 761 7008
rect 421 6916 761 6956
rect 421 1624 550 6916
rect 1374 4490 1498 4530
rect 1374 4438 1410 4490
rect 1462 4438 1498 4490
rect 1374 4272 1498 4438
rect 1374 4220 1410 4272
rect 1462 4220 1498 4272
rect 1374 4180 1498 4220
rect 1635 3830 1760 3869
rect 1635 3774 1670 3830
rect 1726 3774 1760 3830
rect 1635 3653 1760 3774
rect 860 3583 984 3623
rect 860 3531 896 3583
rect 948 3531 984 3583
rect 860 3365 984 3531
rect 1633 3612 1762 3653
rect 1633 3556 1670 3612
rect 1726 3556 1762 3612
rect 1145 3392 1270 3393
rect 860 3313 896 3365
rect 948 3313 984 3365
rect 860 3273 984 3313
rect 1143 3354 1272 3392
rect 1143 3298 1180 3354
rect 1236 3298 1272 3354
rect 421 1572 459 1624
rect 511 1572 550 1624
rect 421 1406 550 1572
rect 421 1359 459 1406
rect 423 1354 459 1359
rect 511 1359 550 1406
rect 1143 3136 1272 3298
rect 1143 3080 1180 3136
rect 1236 3080 1272 3136
rect 1143 1413 1272 3080
rect 1633 1615 1762 3556
rect 511 1354 547 1359
rect 423 1314 547 1354
rect 1143 1280 1762 1413
<< via2 >>
rect 457 8301 513 8303
rect 457 8249 459 8301
rect 459 8249 511 8301
rect 511 8249 513 8301
rect 457 8247 513 8249
rect 664 8301 720 8303
rect 664 8249 666 8301
rect 666 8249 718 8301
rect 718 8249 720 8301
rect 664 8247 720 8249
rect 457 8083 513 8085
rect 457 8031 459 8083
rect 459 8031 511 8083
rect 511 8031 513 8083
rect 457 8029 513 8031
rect 664 8083 720 8085
rect 664 8031 666 8083
rect 666 8031 718 8083
rect 718 8031 720 8083
rect 664 8029 720 8031
rect 457 7865 513 7867
rect 457 7813 459 7865
rect 459 7813 511 7865
rect 511 7813 513 7865
rect 457 7811 513 7813
rect 664 7865 720 7867
rect 664 7813 666 7865
rect 666 7813 718 7865
rect 718 7813 720 7865
rect 664 7811 720 7813
rect 457 7647 513 7649
rect 457 7595 459 7647
rect 459 7595 511 7647
rect 511 7595 513 7647
rect 457 7593 513 7595
rect 664 7647 720 7649
rect 664 7595 666 7647
rect 666 7595 718 7647
rect 718 7595 720 7647
rect 664 7593 720 7595
rect 1184 8278 1240 8280
rect 1184 8226 1186 8278
rect 1186 8226 1238 8278
rect 1238 8226 1240 8278
rect 1184 8224 1240 8226
rect 1184 8060 1240 8062
rect 1184 8008 1186 8060
rect 1186 8008 1238 8060
rect 1238 8008 1240 8060
rect 1184 8006 1240 8008
rect 1184 7842 1240 7844
rect 1184 7790 1186 7842
rect 1186 7790 1238 7842
rect 1238 7790 1240 7842
rect 1184 7788 1240 7790
rect 1184 7624 1240 7626
rect 1184 7572 1186 7624
rect 1186 7572 1238 7624
rect 1238 7572 1240 7624
rect 1184 7570 1240 7572
rect 1670 3774 1726 3830
rect 1670 3556 1726 3612
rect 1180 3298 1236 3354
rect 1180 3080 1236 3136
<< metal3 >>
rect -1 8303 1824 8427
rect -1 8247 457 8303
rect 513 8247 664 8303
rect 720 8280 1824 8303
rect 720 8247 1184 8280
rect -1 8224 1184 8247
rect 1240 8224 1824 8280
rect -1 8085 1824 8224
rect -1 8029 457 8085
rect 513 8029 664 8085
rect 720 8062 1824 8085
rect 720 8029 1184 8062
rect -1 8006 1184 8029
rect 1240 8006 1824 8062
rect -1 7867 1824 8006
rect -1 7811 457 7867
rect 513 7811 664 7867
rect 720 7844 1824 7867
rect 720 7811 1184 7844
rect -1 7788 1184 7811
rect 1240 7788 1824 7844
rect -1 7649 1824 7788
rect -1 7593 457 7649
rect 513 7593 664 7649
rect 720 7626 1824 7649
rect 720 7593 1184 7626
rect -1 7570 1184 7593
rect 1240 7570 1824 7626
rect -1 7519 1824 7570
rect -1 4458 1685 7181
rect 1635 3830 1761 3869
rect 1635 3774 1670 3830
rect 1726 3774 1761 3830
rect 1635 3760 1761 3774
rect 6 3626 1762 3760
rect 1635 3612 1761 3626
rect 1635 3556 1670 3612
rect 1726 3556 1761 3612
rect 1635 3517 1761 3556
rect 1145 3392 1271 3393
rect 15 3354 1815 3392
rect 15 3298 1180 3354
rect 1236 3298 1815 3354
rect 15 3259 1815 3298
rect 1145 3136 1271 3259
rect 1145 3080 1180 3136
rect 1236 3080 1271 3136
rect 1145 3041 1271 3080
use M1_NWELL$$47505452_256x8m81  M1_NWELL$$47505452_256x8m81_0
timestamp 1669390400
transform 1 0 334 0 1 4985
box -221 -1860 221 1860
use M1_POLY2$$46559276_256x8m81_0  M1_POLY2$$46559276_256x8m81_0_0
timestamp 1669390400
transform 1 0 1151 0 1 6982
box 0 0 1 1
use M1_POLY2$$46559276_256x8m81_0  M1_POLY2$$46559276_256x8m81_0_1
timestamp 1669390400
transform 1 0 641 0 1 6982
box 0 0 1 1
use M1_PSUB$$47335468_256x8m81  M1_PSUB$$47335468_256x8m81_0
timestamp 1669390400
transform 1 0 395 0 1 7819
box -79 -572 80 572
use M2_M1$$34864172_256x8m81  M2_M1$$34864172_256x8m81_0
timestamp 1669390400
transform 1 0 591 0 1 6982
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 1489
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1669390400
transform 1 0 922 0 1 3448
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_2
timestamp 1669390400
transform 1 0 1436 0 1 4355
box 0 0 1 1
use M2_M1$$43376684_256x8m81  M2_M1$$43376684_256x8m81_0
timestamp 1669390400
transform 1 0 1219 0 1 5810
box -63 -828 64 828
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 7948
box 0 0 1 1
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_1
timestamp 1669390400
transform 1 0 692 0 1 7948
box 0 0 1 1
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_2
timestamp 1669390400
transform 1 0 1212 0 1 7925
box 0 0 1 1
use M2_M1$$47500332_256x8m81  M2_M1$$47500332_256x8m81_0
timestamp 1669390400
transform 1 0 705 0 1 5584
box -64 -1046 64 1046
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_0
timestamp 1669390400
transform 1 0 1698 0 1 3693
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_1
timestamp 1669390400
transform 1 0 1208 0 1 3217
box 0 0 1 1
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_0
timestamp 1669390400
transform 1 0 485 0 1 7948
box 0 0 1 1
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_1
timestamp 1669390400
transform 1 0 692 0 1 7948
box 0 0 1 1
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_2
timestamp 1669390400
transform 1 0 1212 0 1 7925
box 0 0 1 1
use M3_M2$$47644716_256x8m81  M3_M2$$47644716_256x8m81_0
timestamp 1669390400
transform 1 0 705 0 1 5584
box -65 -1046 65 1046
use M3_M2$$47645740_256x8m81  M3_M2$$47645740_256x8m81_0
timestamp 1669390400
transform 1 0 1219 0 1 5810
box -65 -828 65 828
use alatch_256x8m81  alatch_256x8m81_0
timestamp 1669390400
transform 1 0 70 0 1 -632
box -90 -1 1692 2968
use nmos_1p2$$47502380_256x8m81  nmos_1p2$$47502380_256x8m81_0
timestamp 1669390400
transform 1 0 1296 0 1 7202
box -119 -74 177 1116
use nmos_5p04310590878172_256x8m81  nmos_5p04310590878172_256x8m81_0
timestamp 1669390400
transform 1 0 751 0 1 7123
box -88 -44 208 1452
use pmos_1p2$$47503404_256x8m81  pmos_1p2$$47503404_256x8m81_0
timestamp 1669390400
transform 1 0 782 0 1 3264
box -286 -141 344 3658
use pmos_1p2$$47504428_256x8m81  pmos_1p2$$47504428_256x8m81_0
timestamp 1669390400
transform 1 0 1296 0 1 4171
box -286 -142 343 2752
<< properties >>
string GDS_END 563040
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 560476
<< end >>
