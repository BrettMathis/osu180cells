magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 2998 1094
<< pwell >>
rect -86 -86 2998 453
<< mvnmos >>
rect 168 156 288 314
rect 428 156 548 296
rect 644 156 764 296
rect 812 156 932 296
rect 1036 156 1156 296
rect 1204 156 1324 296
rect 1372 156 1492 296
rect 1632 156 1752 314
rect 1800 156 1920 314
rect 2216 69 2336 333
rect 2440 69 2560 333
rect 2664 69 2784 333
<< mvpmos >>
rect 124 664 244 940
rect 492 740 612 940
rect 804 664 924 864
rect 972 664 1092 864
rect 1196 664 1316 864
rect 1364 664 1484 864
rect 1588 664 1708 864
rect 1848 664 1968 940
rect 2216 574 2336 940
rect 2440 574 2560 940
rect 2664 574 2784 940
<< mvndiff >>
rect 80 215 168 314
rect 80 169 93 215
rect 139 169 168 215
rect 80 156 168 169
rect 288 296 368 314
rect 1552 296 1632 314
rect 288 215 428 296
rect 288 169 317 215
rect 363 169 428 215
rect 288 156 428 169
rect 548 156 644 296
rect 764 156 812 296
rect 932 215 1036 296
rect 932 169 961 215
rect 1007 169 1036 215
rect 932 156 1036 169
rect 1156 156 1204 296
rect 1324 156 1372 296
rect 1492 215 1632 296
rect 1492 169 1521 215
rect 1567 169 1632 215
rect 1492 156 1632 169
rect 1752 156 1800 314
rect 1920 215 2008 314
rect 1920 169 1949 215
rect 1995 169 2008 215
rect 1920 156 2008 169
rect 2128 309 2216 333
rect 2128 169 2141 309
rect 2187 169 2216 309
rect 2128 69 2216 169
rect 2336 295 2440 333
rect 2336 155 2365 295
rect 2411 155 2440 295
rect 2336 69 2440 155
rect 2560 309 2664 333
rect 2560 169 2589 309
rect 2635 169 2664 309
rect 2560 69 2664 169
rect 2784 309 2872 333
rect 2784 169 2813 309
rect 2859 169 2872 309
rect 2784 69 2872 169
<< mvpdiff >>
rect 672 941 744 954
rect 672 940 685 941
rect 36 851 124 940
rect 36 711 49 851
rect 95 711 124 851
rect 36 664 124 711
rect 244 927 332 940
rect 244 787 273 927
rect 319 787 332 927
rect 244 664 332 787
rect 404 833 492 940
rect 404 787 417 833
rect 463 787 492 833
rect 404 740 492 787
rect 612 895 685 940
rect 731 895 744 941
rect 612 864 744 895
rect 1768 864 1848 940
rect 612 740 804 864
rect 724 664 804 740
rect 924 664 972 864
rect 1092 851 1196 864
rect 1092 711 1121 851
rect 1167 711 1196 851
rect 1092 664 1196 711
rect 1316 664 1364 864
rect 1484 851 1588 864
rect 1484 711 1513 851
rect 1559 711 1588 851
rect 1484 664 1588 711
rect 1708 851 1848 864
rect 1708 711 1773 851
rect 1819 711 1848 851
rect 1708 664 1848 711
rect 1968 927 2056 940
rect 1968 787 1997 927
rect 2043 787 2056 927
rect 1968 664 2056 787
rect 2128 851 2216 940
rect 2128 711 2141 851
rect 2187 711 2216 851
rect 2128 574 2216 711
rect 2336 927 2440 940
rect 2336 787 2365 927
rect 2411 787 2440 927
rect 2336 574 2440 787
rect 2560 851 2664 940
rect 2560 711 2589 851
rect 2635 711 2664 851
rect 2560 574 2664 711
rect 2784 927 2872 940
rect 2784 787 2813 927
rect 2859 787 2872 927
rect 2784 574 2872 787
<< mvndiffc >>
rect 93 169 139 215
rect 317 169 363 215
rect 961 169 1007 215
rect 1521 169 1567 215
rect 1949 169 1995 215
rect 2141 169 2187 309
rect 2365 155 2411 295
rect 2589 169 2635 309
rect 2813 169 2859 309
<< mvpdiffc >>
rect 49 711 95 851
rect 273 787 319 927
rect 417 787 463 833
rect 685 895 731 941
rect 1121 711 1167 851
rect 1513 711 1559 851
rect 1773 711 1819 851
rect 1997 787 2043 927
rect 2141 711 2187 851
rect 2365 787 2411 927
rect 2589 711 2635 851
rect 2813 787 2859 927
<< polysilicon >>
rect 124 940 244 984
rect 492 940 612 984
rect 1848 940 1968 984
rect 2216 940 2336 984
rect 2440 940 2560 984
rect 2664 940 2784 984
rect 804 864 924 908
rect 972 864 1092 908
rect 1196 864 1316 908
rect 1364 864 1484 908
rect 1588 864 1708 908
rect 492 696 612 740
rect 124 620 244 664
rect 168 501 244 620
rect 492 514 548 696
rect 804 620 924 664
rect 972 620 1092 664
rect 804 514 844 620
rect 168 455 185 501
rect 231 455 244 501
rect 168 358 244 455
rect 428 501 548 514
rect 428 455 473 501
rect 519 455 548 501
rect 168 314 288 358
rect 428 296 548 455
rect 692 501 844 514
rect 692 455 705 501
rect 751 474 844 501
rect 892 501 964 514
rect 751 455 764 474
rect 692 340 764 455
rect 892 455 905 501
rect 951 455 964 501
rect 892 442 964 455
rect 1012 501 1092 620
rect 1196 620 1316 664
rect 1364 620 1484 664
rect 1196 514 1236 620
rect 1012 455 1025 501
rect 1071 455 1092 501
rect 1012 442 1092 455
rect 1164 501 1236 514
rect 1164 455 1177 501
rect 1223 455 1236 501
rect 1414 508 1484 620
rect 1414 501 1486 508
rect 1414 482 1427 501
rect 1164 442 1236 455
rect 1284 455 1427 482
rect 1473 455 1486 501
rect 1284 442 1486 455
rect 1588 501 1708 664
rect 1588 455 1601 501
rect 1647 455 1708 501
rect 1588 442 1708 455
rect 892 340 932 442
rect 644 296 764 340
rect 812 296 932 340
rect 1036 340 1092 442
rect 1284 340 1324 442
rect 1632 358 1708 442
rect 1848 620 1968 664
rect 1848 501 1920 620
rect 1848 455 1861 501
rect 1907 455 1920 501
rect 1848 358 1920 455
rect 1036 296 1156 340
rect 1204 296 1324 340
rect 1372 296 1492 340
rect 1632 314 1752 358
rect 1800 314 1920 358
rect 2216 530 2336 574
rect 2216 501 2288 530
rect 2440 514 2560 574
rect 2664 514 2784 574
rect 2216 455 2229 501
rect 2275 455 2288 501
rect 2216 377 2288 455
rect 2389 501 2784 514
rect 2389 455 2402 501
rect 2448 455 2784 501
rect 2389 442 2784 455
rect 2216 333 2336 377
rect 2440 333 2560 442
rect 2664 333 2784 442
rect 168 112 288 156
rect 428 112 548 156
rect 644 112 764 156
rect 812 112 932 156
rect 1036 112 1156 156
rect 1204 112 1324 156
rect 429 64 548 112
rect 1372 64 1492 156
rect 1632 112 1752 156
rect 1800 112 1920 156
rect 429 24 1492 64
rect 2216 25 2336 69
rect 2440 25 2560 69
rect 2664 25 2784 69
<< polycontact >>
rect 185 455 231 501
rect 473 455 519 501
rect 705 455 751 501
rect 905 455 951 501
rect 1025 455 1071 501
rect 1177 455 1223 501
rect 1427 455 1473 501
rect 1601 455 1647 501
rect 1861 455 1907 501
rect 2229 455 2275 501
rect 2402 455 2448 501
<< metal1 >>
rect 0 941 2912 1098
rect 0 927 685 941
rect 0 918 273 927
rect 49 851 95 862
rect 319 918 685 927
rect 731 927 2912 941
rect 731 918 1997 927
rect 685 884 731 895
rect 1121 851 1167 862
rect 273 776 319 787
rect 417 838 463 844
rect 417 833 1121 838
rect 463 792 1121 833
rect 417 776 463 787
rect 498 730 1071 746
rect 95 711 1071 730
rect 49 700 1071 711
rect 49 684 533 700
rect 49 215 139 684
rect 185 501 231 512
rect 366 501 530 542
rect 366 455 473 501
rect 519 455 530 501
rect 590 501 642 654
rect 814 501 951 542
rect 590 455 705 501
rect 751 455 762 501
rect 814 455 905 501
rect 185 398 231 455
rect 814 398 951 455
rect 1025 501 1071 700
rect 1121 604 1167 711
rect 1513 851 1559 918
rect 1513 700 1559 711
rect 1773 851 1819 862
rect 2043 918 2365 927
rect 1997 776 2043 787
rect 2141 851 2187 862
rect 1819 711 1999 730
rect 1773 684 1999 711
rect 2411 918 2813 927
rect 2365 776 2411 787
rect 2589 851 2635 862
rect 2187 711 2448 730
rect 2141 684 2448 711
rect 1121 558 1647 604
rect 1025 444 1071 455
rect 1177 501 1223 512
rect 1177 398 1223 455
rect 185 352 1223 398
rect 1269 226 1315 558
rect 1427 501 1473 512
rect 1427 398 1473 455
rect 1601 501 1647 558
rect 1601 444 1647 455
rect 1822 501 1907 542
rect 1822 455 1861 501
rect 1427 352 1642 398
rect 1822 354 1907 455
rect 1953 512 1999 684
rect 1953 501 2275 512
rect 1953 455 2229 501
rect 1953 444 2275 455
rect 2402 501 2448 684
rect 1596 308 1642 352
rect 1953 308 1999 444
rect 2402 398 2448 455
rect 2859 918 2912 927
rect 2813 776 2859 787
rect 2589 430 2635 711
rect 1596 262 1999 308
rect 49 169 93 215
rect 49 158 139 169
rect 317 215 363 226
rect 317 90 363 169
rect 961 215 1315 226
rect 1007 169 1315 215
rect 961 158 1315 169
rect 1521 215 1567 226
rect 1521 90 1567 169
rect 1949 215 1999 262
rect 1995 169 1999 215
rect 1949 158 1999 169
rect 2141 352 2448 398
rect 2141 309 2187 352
rect 2494 309 2635 430
rect 2141 158 2187 169
rect 2365 295 2411 306
rect 2494 242 2589 309
rect 2589 158 2635 169
rect 2813 309 2859 320
rect 2365 90 2411 155
rect 2813 90 2859 169
rect 0 -90 2912 90
<< labels >>
flabel metal1 s 590 501 642 654 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 814 512 951 542 0 FreeSans 200 0 0 0 E
port 2 nsew clock input
flabel metal1 s 2589 430 2635 862 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 366 455 530 542 0 FreeSans 200 0 0 0 RN
port 3 nsew default input
flabel metal1 s 1822 354 1907 542 0 FreeSans 200 0 0 0 SETN
port 4 nsew default input
flabel metal1 s 0 918 2912 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 2813 306 2859 320 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 590 455 762 501 1 D
port 1 nsew default input
rlabel metal1 s 1177 398 1223 512 1 E
port 2 nsew clock input
rlabel metal1 s 814 398 951 512 1 E
port 2 nsew clock input
rlabel metal1 s 185 398 231 512 1 E
port 2 nsew clock input
rlabel metal1 s 185 352 1223 398 1 E
port 2 nsew clock input
rlabel metal1 s 2494 242 2635 430 1 Q
port 5 nsew default output
rlabel metal1 s 2589 158 2635 242 1 Q
port 5 nsew default output
rlabel metal1 s 2813 884 2859 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2365 884 2411 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1997 884 2043 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1513 884 1559 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 685 884 731 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 884 319 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2813 776 2859 884 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2365 776 2411 884 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1997 776 2043 884 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1513 776 1559 884 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 776 319 884 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1513 700 1559 776 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2813 226 2859 306 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2365 226 2411 306 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2813 90 2859 226 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2365 90 2411 226 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1521 90 1567 226 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 317 90 363 226 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2912 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2912 1008
string GDS_END 1019702
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1012292
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
