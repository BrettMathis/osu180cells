VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ffra
  CLASS BLOCK ;
  FOREIGN ffra ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 75.040 900.000 75.600 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 224.560 900.000 225.120 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 374.080 900.000 374.640 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 896.000 523.600 900.000 524.160 ;
    END
  END a[3]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 75.040 4.000 75.600 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 224.560 4.000 225.120 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 374.080 4.000 374.640 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET3 ;
        RECT 0.000 523.600 4.000 524.160 ;
    END
  END b[3]
  PIN ci[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 225.680 0.000 226.240 4.000 ;
    END
  END ci[0]
  PIN ci[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 315.280 0.000 315.840 4.000 ;
    END
  END ci[1]
  PIN ci[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 404.880 0.000 405.440 4.000 ;
    END
  END ci[2]
  PIN ci[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 494.480 0.000 495.040 4.000 ;
    END
  END ci[3]
  PIN ci[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 584.080 0.000 584.640 4.000 ;
    END
  END ci[4]
  PIN ci[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 673.680 0.000 674.240 4.000 ;
    END
  END ci[5]
  PIN ci[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 763.280 0.000 763.840 4.000 ;
    END
  END ci[6]
  PIN ci[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 852.880 0.000 853.440 4.000 ;
    END
  END ci[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 46.480 0.000 47.040 4.000 ;
    END
  END clk
  PIN o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 57.680 596.000 58.240 600.000 ;
    END
  END o[0]
  PIN o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 169.680 596.000 170.240 600.000 ;
    END
  END o[1]
  PIN o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 281.680 596.000 282.240 600.000 ;
    END
  END o[2]
  PIN o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 393.680 596.000 394.240 600.000 ;
    END
  END o[3]
  PIN o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 505.680 596.000 506.240 600.000 ;
    END
  END o[4]
  PIN o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 617.680 596.000 618.240 600.000 ;
    END
  END o[5]
  PIN o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 729.680 596.000 730.240 600.000 ;
    END
  END o[6]
  PIN o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 841.680 596.000 842.240 600.000 ;
    END
  END o[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 136.080 0.000 136.640 4.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET4 ;
        RECT 16.720 24.300 18.320 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 170.320 24.300 171.920 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 323.920 24.300 325.520 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 477.520 24.300 479.120 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 631.120 24.300 632.720 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 784.720 24.300 786.320 572.250 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET4 ;
        RECT 93.520 24.300 95.120 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 247.120 24.300 248.720 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 400.720 24.300 402.320 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 554.320 24.300 555.920 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 707.920 24.300 709.520 572.250 ;
    END
    PORT
      LAYER MET4 ;
        RECT 861.520 24.300 863.120 572.250 ;
    END
  END vss
  OBS
      LAYER MET1 ;
        RECT 1.200 24.300 898.800 572.250 ;
      LAYER MET2 ;
        RECT 3.360 595.700 57.380 596.820 ;
        RECT 58.540 595.700 169.380 596.820 ;
        RECT 170.540 595.700 281.380 596.820 ;
        RECT 282.540 595.700 393.380 596.820 ;
        RECT 394.540 595.700 505.380 596.820 ;
        RECT 506.540 595.700 617.380 596.820 ;
        RECT 618.540 595.700 729.380 596.820 ;
        RECT 730.540 595.700 841.380 596.820 ;
        RECT 842.540 595.700 897.590 596.820 ;
        RECT 3.360 4.300 897.590 595.700 ;
        RECT 3.360 4.000 46.180 4.300 ;
        RECT 47.340 4.000 135.780 4.300 ;
        RECT 136.940 4.000 225.380 4.300 ;
        RECT 226.540 4.000 314.980 4.300 ;
        RECT 316.140 4.000 404.580 4.300 ;
        RECT 405.740 4.000 494.180 4.300 ;
        RECT 495.340 4.000 583.780 4.300 ;
        RECT 584.940 4.000 673.380 4.300 ;
        RECT 674.540 4.000 762.980 4.300 ;
        RECT 764.140 4.000 852.580 4.300 ;
        RECT 853.740 4.000 897.590 4.300 ;
      LAYER MET3 ;
        RECT 3.450 524.460 897.590 572.090 ;
        RECT 4.300 523.300 895.700 524.460 ;
        RECT 3.450 374.940 897.590 523.300 ;
        RECT 4.300 373.780 895.700 374.940 ;
        RECT 3.450 225.420 897.590 373.780 ;
        RECT 4.300 224.260 895.700 225.420 ;
        RECT 3.450 75.900 897.590 224.260 ;
        RECT 4.300 74.740 895.700 75.900 ;
        RECT 3.450 24.460 897.590 74.740 ;
      LAYER MET4 ;
        RECT 332.780 146.810 400.420 286.070 ;
        RECT 402.620 146.810 477.220 286.070 ;
        RECT 479.420 146.810 554.020 286.070 ;
        RECT 556.220 146.810 588.980 286.070 ;
  END
END ffra
END LIBRARY

