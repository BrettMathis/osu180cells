magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 5798 1094
<< pwell >>
rect -86 -86 5798 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
rect 1468 69 1588 333
rect 1692 69 1812 333
rect 1916 69 2036 333
rect 2140 69 2260 333
rect 2364 69 2484 333
rect 2588 69 2708 333
rect 2916 69 3036 333
rect 3140 69 3260 333
rect 3364 69 3484 333
rect 3588 69 3708 333
rect 3812 69 3932 333
rect 4036 69 4156 333
rect 4260 69 4380 333
rect 4484 69 4604 333
rect 4708 69 4828 333
rect 4932 69 5052 333
rect 5156 69 5276 333
rect 5380 69 5500 333
<< mvpmos >>
rect 134 573 234 939
rect 348 573 448 939
rect 582 573 682 939
rect 806 573 906 939
rect 1030 573 1130 939
rect 1244 573 1344 939
rect 1478 573 1578 939
rect 1702 573 1802 939
rect 1926 573 2026 939
rect 2140 573 2240 939
rect 2384 573 2484 939
rect 2588 573 2688 939
rect 2936 573 3036 939
rect 3160 573 3260 939
rect 3374 573 3474 939
rect 3598 573 3698 939
rect 3822 573 3922 939
rect 4046 573 4146 939
rect 4280 573 4380 939
rect 4494 573 4594 939
rect 4718 573 4818 939
rect 4942 573 5042 939
rect 5166 573 5266 939
rect 5380 573 5480 939
<< mvndiff >>
rect 36 297 124 333
rect 36 157 49 297
rect 95 157 124 297
rect 36 69 124 157
rect 244 203 348 333
rect 244 157 273 203
rect 319 157 348 203
rect 244 69 348 157
rect 468 297 572 333
rect 468 157 497 297
rect 543 157 572 297
rect 468 69 572 157
rect 692 203 796 333
rect 692 157 721 203
rect 767 157 796 203
rect 692 69 796 157
rect 916 297 1020 333
rect 916 157 945 297
rect 991 157 1020 297
rect 916 69 1020 157
rect 1140 203 1244 333
rect 1140 157 1169 203
rect 1215 157 1244 203
rect 1140 69 1244 157
rect 1364 297 1468 333
rect 1364 157 1393 297
rect 1439 157 1468 297
rect 1364 69 1468 157
rect 1588 203 1692 333
rect 1588 157 1617 203
rect 1663 157 1692 203
rect 1588 69 1692 157
rect 1812 297 1916 333
rect 1812 157 1841 297
rect 1887 157 1916 297
rect 1812 69 1916 157
rect 2036 203 2140 333
rect 2036 157 2065 203
rect 2111 157 2140 203
rect 2036 69 2140 157
rect 2260 297 2364 333
rect 2260 157 2289 297
rect 2335 157 2364 297
rect 2260 69 2364 157
rect 2484 203 2588 333
rect 2484 157 2513 203
rect 2559 157 2588 203
rect 2484 69 2588 157
rect 2708 203 2916 333
rect 2708 157 2841 203
rect 2887 157 2916 203
rect 2708 69 2916 157
rect 3036 306 3140 333
rect 3036 260 3065 306
rect 3111 260 3140 306
rect 3036 69 3140 260
rect 3260 203 3364 333
rect 3260 157 3289 203
rect 3335 157 3364 203
rect 3260 69 3364 157
rect 3484 274 3588 333
rect 3484 228 3513 274
rect 3559 228 3588 274
rect 3484 69 3588 228
rect 3708 203 3812 333
rect 3708 157 3737 203
rect 3783 157 3812 203
rect 3708 69 3812 157
rect 3932 274 4036 333
rect 3932 228 3961 274
rect 4007 228 4036 274
rect 3932 69 4036 228
rect 4156 203 4260 333
rect 4156 157 4185 203
rect 4231 157 4260 203
rect 4156 69 4260 157
rect 4380 274 4484 333
rect 4380 228 4409 274
rect 4455 228 4484 274
rect 4380 69 4484 228
rect 4604 203 4708 333
rect 4604 157 4633 203
rect 4679 157 4708 203
rect 4604 69 4708 157
rect 4828 274 4932 333
rect 4828 228 4857 274
rect 4903 228 4932 274
rect 4828 69 4932 228
rect 5052 203 5156 333
rect 5052 157 5081 203
rect 5127 157 5156 203
rect 5052 69 5156 157
rect 5276 306 5380 333
rect 5276 260 5305 306
rect 5351 260 5380 306
rect 5276 69 5380 260
rect 5500 203 5588 333
rect 5500 157 5529 203
rect 5575 157 5588 203
rect 5500 69 5588 157
<< mvpdiff >>
rect 46 775 134 939
rect 46 635 59 775
rect 105 635 134 775
rect 46 573 134 635
rect 234 573 348 939
rect 448 867 582 939
rect 448 727 477 867
rect 523 727 582 867
rect 448 573 582 727
rect 682 573 806 939
rect 906 775 1030 939
rect 906 635 935 775
rect 981 635 1030 775
rect 906 573 1030 635
rect 1130 573 1244 939
rect 1344 867 1478 939
rect 1344 727 1373 867
rect 1419 727 1478 867
rect 1344 573 1478 727
rect 1578 573 1702 939
rect 1802 573 1926 939
rect 2026 755 2140 939
rect 2026 615 2065 755
rect 2111 615 2140 755
rect 2026 573 2140 615
rect 2240 847 2384 939
rect 2240 707 2269 847
rect 2315 707 2384 847
rect 2240 573 2384 707
rect 2484 755 2588 939
rect 2484 615 2513 755
rect 2559 615 2588 755
rect 2484 573 2588 615
rect 2688 858 2776 939
rect 2688 812 2717 858
rect 2763 812 2776 858
rect 2688 573 2776 812
rect 2848 753 2936 939
rect 2848 707 2861 753
rect 2907 707 2936 753
rect 2848 573 2936 707
rect 3036 681 3160 939
rect 3036 635 3065 681
rect 3111 635 3160 681
rect 3036 573 3160 635
rect 3260 753 3374 939
rect 3260 707 3289 753
rect 3335 707 3374 753
rect 3260 573 3374 707
rect 3474 681 3598 939
rect 3474 635 3503 681
rect 3549 635 3598 681
rect 3474 573 3598 635
rect 3698 573 3822 939
rect 3922 573 4046 939
rect 4146 887 4280 939
rect 4146 841 4175 887
rect 4221 841 4280 887
rect 4146 573 4280 841
rect 4380 573 4494 939
rect 4594 740 4718 939
rect 4594 694 4623 740
rect 4669 694 4718 740
rect 4594 573 4718 694
rect 4818 573 4942 939
rect 5042 926 5166 939
rect 5042 786 5071 926
rect 5117 786 5166 926
rect 5042 573 5166 786
rect 5266 573 5380 939
rect 5480 834 5568 939
rect 5480 694 5509 834
rect 5555 694 5568 834
rect 5480 573 5568 694
<< mvndiffc >>
rect 49 157 95 297
rect 273 157 319 203
rect 497 157 543 297
rect 721 157 767 203
rect 945 157 991 297
rect 1169 157 1215 203
rect 1393 157 1439 297
rect 1617 157 1663 203
rect 1841 157 1887 297
rect 2065 157 2111 203
rect 2289 157 2335 297
rect 2513 157 2559 203
rect 2841 157 2887 203
rect 3065 260 3111 306
rect 3289 157 3335 203
rect 3513 228 3559 274
rect 3737 157 3783 203
rect 3961 228 4007 274
rect 4185 157 4231 203
rect 4409 228 4455 274
rect 4633 157 4679 203
rect 4857 228 4903 274
rect 5081 157 5127 203
rect 5305 260 5351 306
rect 5529 157 5575 203
<< mvpdiffc >>
rect 59 635 105 775
rect 477 727 523 867
rect 935 635 981 775
rect 1373 727 1419 867
rect 2065 615 2111 755
rect 2269 707 2315 847
rect 2513 615 2559 755
rect 2717 812 2763 858
rect 2861 707 2907 753
rect 3065 635 3111 681
rect 3289 707 3335 753
rect 3503 635 3549 681
rect 4175 841 4221 887
rect 4623 694 4669 740
rect 5071 786 5117 926
rect 5509 694 5555 834
<< polysilicon >>
rect 134 939 234 983
rect 348 939 448 983
rect 582 939 682 983
rect 806 939 906 983
rect 1030 939 1130 983
rect 1244 939 1344 983
rect 1478 939 1578 983
rect 1702 939 1802 983
rect 1926 939 2026 983
rect 2140 939 2240 983
rect 2384 939 2484 983
rect 2588 939 2688 983
rect 2936 939 3036 983
rect 3160 939 3260 983
rect 3374 939 3474 983
rect 3598 939 3698 983
rect 3822 939 3922 983
rect 4046 939 4146 983
rect 4280 939 4380 983
rect 4494 939 4594 983
rect 4718 939 4818 983
rect 4942 939 5042 983
rect 5166 939 5266 983
rect 5380 939 5480 983
rect 134 484 234 573
rect 134 438 175 484
rect 221 438 234 484
rect 134 377 234 438
rect 348 513 448 573
rect 582 513 682 573
rect 348 484 682 513
rect 348 438 377 484
rect 423 441 682 484
rect 423 438 468 441
rect 124 333 244 377
rect 348 333 468 438
rect 572 377 682 441
rect 806 513 906 573
rect 1030 513 1130 573
rect 806 500 1130 513
rect 806 454 819 500
rect 865 454 1130 500
rect 806 441 1130 454
rect 806 377 916 441
rect 572 333 692 377
rect 796 333 916 377
rect 1020 377 1130 441
rect 1244 513 1344 573
rect 1478 513 1578 573
rect 1244 484 1578 513
rect 1244 438 1257 484
rect 1303 441 1578 484
rect 1303 438 1364 441
rect 1020 333 1140 377
rect 1244 333 1364 438
rect 1468 377 1578 441
rect 1702 500 1802 573
rect 1702 454 1715 500
rect 1761 454 1802 500
rect 1702 377 1802 454
rect 1926 513 2026 573
rect 2140 513 2240 573
rect 1926 500 2240 513
rect 1926 454 2065 500
rect 2111 497 2240 500
rect 2384 513 2484 573
rect 2588 513 2688 573
rect 2384 500 2688 513
rect 2384 497 2513 500
rect 2111 484 2513 497
rect 2111 454 2289 484
rect 1926 441 2289 454
rect 1926 377 2036 441
rect 1468 333 1588 377
rect 1692 333 1812 377
rect 1916 333 2036 377
rect 2140 438 2289 441
rect 2335 454 2513 484
rect 2559 454 2688 500
rect 2335 441 2688 454
rect 2335 438 2484 441
rect 2140 425 2484 438
rect 2140 333 2260 425
rect 2364 333 2484 425
rect 2588 377 2688 441
rect 2936 513 3036 573
rect 3160 513 3260 573
rect 3374 513 3474 573
rect 2936 500 3474 513
rect 2936 454 3065 500
rect 3111 454 3289 500
rect 3335 497 3474 500
rect 3598 497 3698 573
rect 3335 484 3698 497
rect 3335 454 3513 484
rect 2936 441 3513 454
rect 2936 377 3036 441
rect 2588 333 2708 377
rect 2916 333 3036 377
rect 3140 333 3260 441
rect 3364 438 3513 441
rect 3559 438 3698 484
rect 3364 425 3698 438
rect 3364 333 3484 425
rect 3588 377 3698 425
rect 3822 500 3922 573
rect 3822 454 3835 500
rect 3881 454 3922 500
rect 3822 377 3922 454
rect 4046 513 4146 573
rect 4280 513 4380 573
rect 4046 453 4380 513
rect 4046 407 4059 453
rect 4105 441 4380 453
rect 4105 407 4156 441
rect 4046 377 4156 407
rect 3588 333 3708 377
rect 3812 333 3932 377
rect 4036 333 4156 377
rect 4260 333 4380 441
rect 4494 513 4594 573
rect 4718 513 4818 573
rect 4494 500 4818 513
rect 4494 454 4507 500
rect 4553 454 4818 500
rect 4494 441 4818 454
rect 4494 377 4604 441
rect 4484 333 4604 377
rect 4708 377 4818 441
rect 4942 513 5042 573
rect 5166 513 5266 573
rect 4942 453 5266 513
rect 4942 407 4955 453
rect 5001 441 5266 453
rect 5001 407 5052 441
rect 4942 377 5052 407
rect 4708 333 4828 377
rect 4932 333 5052 377
rect 5156 377 5266 441
rect 5380 500 5480 573
rect 5380 454 5393 500
rect 5439 454 5480 500
rect 5380 377 5480 454
rect 5156 333 5276 377
rect 5380 333 5500 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1468 25 1588 69
rect 1692 25 1812 69
rect 1916 25 2036 69
rect 2140 25 2260 69
rect 2364 25 2484 69
rect 2588 25 2708 69
rect 2916 25 3036 69
rect 3140 25 3260 69
rect 3364 25 3484 69
rect 3588 25 3708 69
rect 3812 25 3932 69
rect 4036 25 4156 69
rect 4260 25 4380 69
rect 4484 25 4604 69
rect 4708 25 4828 69
rect 4932 25 5052 69
rect 5156 25 5276 69
rect 5380 25 5500 69
<< polycontact >>
rect 175 438 221 484
rect 377 438 423 484
rect 819 454 865 500
rect 1257 438 1303 484
rect 1715 454 1761 500
rect 2065 454 2111 500
rect 2289 438 2335 484
rect 2513 454 2559 500
rect 3065 454 3111 500
rect 3289 454 3335 500
rect 3513 438 3559 484
rect 3835 454 3881 500
rect 4059 407 4105 453
rect 4507 454 4553 500
rect 4955 407 5001 453
rect 5393 454 5439 500
<< metal1 >>
rect 0 926 5712 1098
rect 0 918 5071 926
rect 477 867 523 918
rect 59 775 105 786
rect 1373 867 1419 918
rect 477 716 523 727
rect 935 775 981 786
rect 105 635 935 670
rect 4175 887 4221 918
rect 1373 716 1419 727
rect 1465 847 2717 858
rect 1465 812 2269 847
rect 1465 670 1511 812
rect 981 635 1511 670
rect 59 624 1511 635
rect 2065 755 2111 766
rect 2315 812 2717 847
rect 2763 812 2774 858
rect 4175 830 4221 841
rect 5117 918 5712 926
rect 2269 696 2315 707
rect 2513 755 2770 766
rect 2111 615 2513 637
rect 2559 637 2770 755
rect 2861 753 4669 784
rect 5071 775 5117 786
rect 5509 834 5555 845
rect 2907 738 3289 753
rect 2861 696 2907 707
rect 3335 740 4669 753
rect 3335 738 4623 740
rect 3289 696 3335 707
rect 4669 694 5509 729
rect 3065 681 3111 692
rect 2559 635 3065 637
rect 3503 681 3549 692
rect 4623 683 5555 694
rect 3111 635 3503 637
rect 3549 635 5531 637
rect 2559 615 5531 635
rect 2065 591 5531 615
rect 164 530 1406 576
rect 164 484 232 530
rect 808 500 876 530
rect 164 438 175 484
rect 221 438 232 484
rect 366 438 377 484
rect 423 438 434 484
rect 808 454 819 500
rect 865 454 876 500
rect 1360 500 1406 530
rect 2065 500 2559 542
rect 366 400 434 438
rect 922 438 1257 484
rect 1303 438 1314 484
rect 1360 454 1715 500
rect 1761 454 1772 500
rect 2111 484 2513 500
rect 2111 454 2289 484
rect 2065 438 2289 454
rect 2335 454 2513 484
rect 2335 438 2559 454
rect 3065 500 3570 542
rect 3111 454 3289 500
rect 3335 484 3570 500
rect 3335 454 3513 484
rect 3065 438 3513 454
rect 3559 438 3570 484
rect 3824 500 5439 545
rect 3824 454 3835 500
rect 3881 499 4507 500
rect 3881 454 3892 499
rect 4398 454 4507 499
rect 4553 499 5393 500
rect 4553 454 4564 499
rect 922 400 968 438
rect 366 354 968 400
rect 3938 407 4059 453
rect 4105 408 4116 453
rect 4944 408 4955 453
rect 4105 407 4955 408
rect 5001 407 5012 453
rect 5393 443 5439 454
rect 3938 362 5012 407
rect 49 297 2886 308
rect 5485 306 5531 591
rect 95 262 497 297
rect 49 146 95 157
rect 273 203 319 214
rect 273 90 319 157
rect 543 262 945 297
rect 497 146 543 157
rect 721 203 767 214
rect 721 90 767 157
rect 991 262 1393 297
rect 945 146 991 157
rect 1169 203 1215 214
rect 1169 90 1215 157
rect 1439 262 1841 297
rect 1393 146 1439 157
rect 1617 203 1663 214
rect 1617 90 1663 157
rect 1887 262 2289 297
rect 1841 146 1887 157
rect 2065 203 2111 214
rect 2065 90 2111 157
rect 2335 262 2886 297
rect 2840 214 2886 262
rect 3054 260 3065 306
rect 3111 274 5305 306
rect 3111 260 3513 274
rect 3502 228 3513 260
rect 3559 260 3961 274
rect 3559 228 3570 260
rect 3950 228 3961 260
rect 4007 260 4409 274
rect 4007 228 4018 260
rect 4398 228 4409 260
rect 4455 260 4857 274
rect 4455 228 4466 260
rect 4846 228 4857 260
rect 4903 260 5305 274
rect 5351 260 5531 306
rect 4903 228 4914 260
rect 2289 146 2335 157
rect 2513 203 2559 214
rect 2513 90 2559 157
rect 2840 203 3335 214
rect 5081 203 5575 214
rect 2840 157 2841 203
rect 2887 157 3289 203
rect 3726 182 3737 203
rect 3335 157 3737 182
rect 3783 182 3794 203
rect 4174 182 4185 203
rect 3783 157 4185 182
rect 4231 182 4242 203
rect 4622 182 4633 203
rect 4231 157 4633 182
rect 4679 182 4690 203
rect 4679 157 5081 182
rect 5127 157 5529 203
rect 2840 136 5575 157
rect 0 -90 5712 90
<< labels >>
flabel metal1 s 3065 438 3570 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 3824 499 5439 545 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 4944 408 5012 453 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 2065 438 2559 542 0 FreeSans 200 0 0 0 B1
port 4 nsew default input
flabel metal1 s 164 530 1406 576 0 FreeSans 200 0 0 0 B2
port 5 nsew default input
flabel metal1 s 922 438 1314 484 0 FreeSans 200 0 0 0 B3
port 6 nsew default input
flabel metal1 s 0 918 5712 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 2513 90 2559 214 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 2513 692 2770 766 0 FreeSans 200 0 0 0 ZN
port 7 nsew default output
rlabel metal1 s 5393 454 5439 499 1 A2
port 2 nsew default input
rlabel metal1 s 4398 454 4564 499 1 A2
port 2 nsew default input
rlabel metal1 s 3824 454 3892 499 1 A2
port 2 nsew default input
rlabel metal1 s 5393 443 5439 454 1 A2
port 2 nsew default input
rlabel metal1 s 3938 408 4116 453 1 A3
port 3 nsew default input
rlabel metal1 s 3938 362 5012 408 1 A3
port 3 nsew default input
rlabel metal1 s 1360 500 1406 530 1 B2
port 5 nsew default input
rlabel metal1 s 808 500 876 530 1 B2
port 5 nsew default input
rlabel metal1 s 164 500 232 530 1 B2
port 5 nsew default input
rlabel metal1 s 1360 454 1772 500 1 B2
port 5 nsew default input
rlabel metal1 s 808 454 876 500 1 B2
port 5 nsew default input
rlabel metal1 s 164 454 232 500 1 B2
port 5 nsew default input
rlabel metal1 s 164 438 232 454 1 B2
port 5 nsew default input
rlabel metal1 s 366 438 434 484 1 B3
port 6 nsew default input
rlabel metal1 s 922 400 968 438 1 B3
port 6 nsew default input
rlabel metal1 s 366 400 434 438 1 B3
port 6 nsew default input
rlabel metal1 s 366 354 968 400 1 B3
port 6 nsew default input
rlabel metal1 s 2065 692 2111 766 1 ZN
port 7 nsew default output
rlabel metal1 s 3503 637 3549 692 1 ZN
port 7 nsew default output
rlabel metal1 s 3065 637 3111 692 1 ZN
port 7 nsew default output
rlabel metal1 s 2513 637 2770 692 1 ZN
port 7 nsew default output
rlabel metal1 s 2065 637 2111 692 1 ZN
port 7 nsew default output
rlabel metal1 s 2065 591 5531 637 1 ZN
port 7 nsew default output
rlabel metal1 s 5485 306 5531 591 1 ZN
port 7 nsew default output
rlabel metal1 s 3054 260 5531 306 1 ZN
port 7 nsew default output
rlabel metal1 s 4846 228 4914 260 1 ZN
port 7 nsew default output
rlabel metal1 s 4398 228 4466 260 1 ZN
port 7 nsew default output
rlabel metal1 s 3950 228 4018 260 1 ZN
port 7 nsew default output
rlabel metal1 s 3502 228 3570 260 1 ZN
port 7 nsew default output
rlabel metal1 s 5071 830 5117 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4175 830 4221 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1373 830 1419 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 477 830 523 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5071 775 5117 830 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1373 775 1419 830 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 477 775 523 830 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1373 716 1419 775 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 477 716 523 775 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2065 90 2111 214 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1617 90 1663 214 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1169 90 1215 214 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 721 90 767 214 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 214 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5712 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5712 1008
string GDS_END 198800
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 188676
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
