magic
tech gf180mcuA
magscale 1 10
timestamp 1669390400
<< psubdiff >>
rect -42 31323 842 31342
rect -42 -23 -23 31323
rect 823 -23 842 31323
rect -42 -42 842 -23
<< psubdiffcont >>
rect -23 -23 823 31323
<< metal1 >>
rect -34 31323 834 31334
rect -34 -23 -23 31323
rect 823 -23 834 31323
rect -34 -34 834 -23
<< properties >>
string GDS_END 1593652
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1412592
<< end >>
