# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__addf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 16.8 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.265 2.33 3.455 2.33 3.455 2.71 2.265 2.71  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.525 2.265 13.85 2.265 13.85 2.71 13.525 2.71  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.547 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.89 2.115 7.975 2.115 11.91 2.115 11.91 1.77 12.11 1.77 12.17 1.77 12.17 2.115 12.55 2.115 12.55 2.345 12.11 2.345 7.975 2.345 3.89 2.345  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.83 2.89 16.145 2.89 16.145 0.845 16.475 0.845 16.475 3.685 15.83 3.685  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.3244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 0.845 0.575 0.845 0.575 3.83 0.15 3.83  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.875 1.595 3.875 1.595 4.59 4.615 4.59 6.625 4.59 6.625 3.61 6.855 3.61 6.855 4.59 7.93 4.59 8.665 4.59 8.665 3.14 8.895 3.14 8.895 4.59 10.705 4.59 10.705 3.505 10.935 3.505 10.935 4.59 11.955 4.59 15.125 4.59 15.125 3.875 15.355 3.875 15.355 4.59 15.795 4.59 16.8 4.59 16.8 5.49 15.795 5.49 11.955 5.49 7.93 5.49 4.615 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 16.8 -0.45 16.8 0.45 15.355 0.45 15.355 1.165 15.125 1.165 15.125 0.45 10.935 0.45 10.935 1.425 10.705 1.425 10.705 0.45 9.095 0.45 9.095 1.425 8.865 1.425 8.865 0.45 6.855 0.45 6.855 1.425 6.625 1.425 6.625 0.45 1.595 0.45 1.595 1.305 1.365 1.305 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.035 2.94 4.615 2.94 4.615 3.79 4.385 3.79 4.385 3.17 1.805 3.17 1.805 2.06 0.87 2.06 0.87 1.655 4.385 1.655 4.385 1.315 4.615 1.315 4.615 1.885 2.035 1.885  ;
        POLYGON 5.605 3.035 7.93 3.035 7.93 3.265 5.835 3.265 5.835 3.845 5.605 3.845  ;
        POLYGON 5.505 1.315 5.735 1.315 5.735 1.655 7.745 1.655 7.745 1.315 7.975 1.315 7.975 1.885 5.505 1.885  ;
        POLYGON 9.685 3.035 11.955 3.035 11.955 3.845 11.725 3.845 11.725 3.265 9.915 3.265 9.915 3.845 9.685 3.845  ;
        POLYGON 9.585 1.315 9.815 1.315 9.815 1.655 11.45 1.655 11.45 1.31 12.11 1.31 12.11 1.54 11.68 1.54 11.68 1.885 9.585 1.885  ;
        POLYGON 5.01 2.575 13.075 2.575 13.075 2.94 14.08 2.94 14.08 2.005 12.945 2.005 12.945 1.315 13.175 1.315 13.175 1.775 15.795 1.775 15.795 2.115 14.31 2.115 14.31 3.17 13.075 3.17 13.075 3.685 12.845 3.685 12.845 2.805 5.01 2.805  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.7 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.425 2.33 4.605 2.33 4.605 2.71 3.425 2.71  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.7 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 2.15 16.11 2.15 16.11 2.71 14.71 2.71  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.525 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.05 1.92 5.83 1.92 9.135 1.92 13.215 1.92 13.59 1.92 13.59 1.77 13.85 1.77 13.85 2.15 13.215 2.15 9.135 2.15 5.83 2.15 5.05 2.15  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.165 0.845 17.77 0.845 17.77 2.71 17.395 2.71 17.395 3.685 17.165 3.685  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 0.845 1.855 0.845 1.855 3.83 1.27 3.83  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.605 4.59 0.605 3.845 0.835 3.845 0.835 4.59 2.645 4.59 2.645 3.845 2.875 3.845 2.875 4.59 5.83 4.59 7.785 4.59 7.785 3.905 8.015 3.905 8.015 4.59 9.035 4.59 10.025 4.59 10.025 3.435 10.255 3.435 10.255 4.59 11.765 4.59 11.765 3.435 11.995 3.435 11.995 4.59 13.115 4.59 15.965 4.59 15.965 3.905 16.195 3.905 16.195 4.59 16.935 4.59 18.185 4.59 18.185 3.845 18.415 3.845 18.415 4.59 19.04 4.59 19.04 5.49 16.935 5.49 13.115 5.49 9.035 5.49 5.83 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 18.735 0.45 18.735 1.165 18.505 1.165 18.505 0.45 16.495 0.45 16.495 1.195 16.265 1.195 16.265 0.45 12.095 0.45 12.095 1.215 11.865 1.215 11.865 0.45 10.255 0.45 10.255 1.215 10.025 1.215 10.025 0.45 8.015 0.45 8.015 1.215 7.785 1.215 7.785 0.45 2.755 0.45 2.755 1.165 2.525 1.165 2.525 0.45 0.515 0.45 0.515 1.165 0.285 1.165 0.285 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.085 1.775 2.965 1.775 2.965 1.37 5.83 1.37 5.83 1.6 3.195 1.6 3.195 2.94 5.545 2.94 5.545 2.875 5.775 2.875 5.775 3.685 5.545 3.685 5.545 3.17 2.965 3.17 2.965 2.115 2.085 2.115  ;
        POLYGON 6.71 2.93 9.035 2.93 9.035 3.74 8.805 3.74 8.805 3.16 6.71 3.16  ;
        POLYGON 6.665 1.315 6.895 1.315 6.895 1.445 8.905 1.445 8.905 1.315 9.135 1.315 9.135 1.675 6.665 1.675  ;
        POLYGON 10.745 2.93 13.115 2.93 13.115 3.74 12.885 3.74 12.885 3.16 10.975 3.16 10.975 3.74 10.745 3.74  ;
        POLYGON 10.745 1.315 10.975 1.315 10.975 1.445 12.985 1.445 12.985 1.315 13.215 1.315 13.215 1.675 10.745 1.675  ;
        POLYGON 6.07 2.47 14.335 2.47 14.335 2.985 16.705 2.985 16.705 1.655 14.05 1.655 14.05 1.37 14.39 1.37 14.39 1.425 16.935 1.425 16.935 3.215 14.105 3.215 14.105 2.7 6.07 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.7 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.705 1.86 6.785 1.86 6.785 2.71 5.705 2.71  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.7 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.965 2.33 18.53 2.33 18.53 2.71 16.965 2.71  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.525 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.33 1.92 8.11 1.92 11.415 1.92 11.91 1.92 11.91 1.77 12.17 1.77 12.17 1.92 15.495 1.92 15.99 1.92 15.99 2.15 15.495 2.15 11.415 2.15 8.11 2.15 7.33 2.15  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.635 2.875 20.725 2.875 20.725 1.655 19.685 1.655 19.685 0.845 19.915 0.845 19.915 1.425 21.925 1.425 21.925 0.845 22.155 0.845 22.155 1.655 21.185 1.655 21.185 2.875 22.105 2.875 22.105 3.685 21.875 3.685 21.875 3.105 19.865 3.105 19.865 3.685 19.635 3.685  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.81585 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.84 2.875 4.015 2.875 4.015 3.685 3.785 3.685 3.785 3.105 1.675 3.105 1.675 3.685 1.445 3.685 1.445 2.875 2.38 2.875 2.38 1.655 1.445 1.655 1.445 0.845 1.675 0.845 1.675 1.425 3.685 1.425 3.685 0.845 3.915 0.845 3.915 1.655 2.84 1.655  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.325 4.59 0.325 3.875 0.555 3.875 0.555 4.59 2.555 4.59 2.555 3.875 2.785 3.875 2.785 4.59 4.905 4.59 4.905 3.875 5.135 3.875 5.135 4.59 8.11 4.59 10.065 4.59 10.065 3.905 10.295 3.905 10.295 4.59 11.37 4.59 12.205 4.59 12.205 3.435 12.435 3.435 12.435 4.59 14.145 4.59 14.145 3.435 14.375 3.435 14.375 4.59 15.395 4.59 18.465 4.59 18.465 3.875 18.695 3.875 18.695 4.59 19.235 4.59 20.75 4.59 20.75 3.875 20.98 3.875 20.98 4.59 22.945 4.59 22.945 3.875 23.175 3.875 23.175 4.59 23.52 4.59 23.52 5.49 19.235 5.49 15.395 5.49 11.37 5.49 8.11 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 23.275 0.45 23.275 1.165 23.045 1.165 23.045 0.45 21.035 0.45 21.035 1.165 20.805 1.165 20.805 0.45 18.795 0.45 18.795 1.165 18.565 1.165 18.565 0.45 14.375 0.45 14.375 1.215 14.145 1.215 14.145 0.45 12.535 0.45 12.535 1.215 12.305 1.215 12.305 0.45 10.295 0.45 10.295 1.215 10.065 1.215 10.065 0.45 5.035 0.45 5.035 1.165 4.805 1.165 4.805 0.45 2.795 0.45 2.795 1.165 2.565 1.165 2.565 0.45 0.555 0.45 0.555 1.165 0.325 1.165 0.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.31 1.83 5.245 1.83 5.245 1.315 8.11 1.315 8.11 1.545 5.475 1.545 5.475 2.94 7.825 2.94 7.825 2.875 8.055 2.875 8.055 3.685 7.825 3.685 7.825 3.17 5.245 3.17 5.245 2.06 4.595 2.06 4.595 2.585 4.31 2.585  ;
        POLYGON 9.045 2.93 11.37 2.93 11.37 3.16 9.275 3.16 9.275 3.74 9.045 3.74  ;
        POLYGON 8.945 1.315 9.175 1.315 9.175 1.445 11.185 1.445 11.185 1.315 11.415 1.315 11.415 1.675 8.945 1.675  ;
        POLYGON 13.125 2.93 15.395 2.93 15.395 3.74 15.165 3.74 15.165 3.16 13.355 3.16 13.355 3.74 13.125 3.74  ;
        POLYGON 13.025 1.315 13.255 1.315 13.255 1.445 15.265 1.445 15.265 1.315 15.495 1.315 15.495 1.675 13.025 1.675  ;
        POLYGON 8.45 2.47 15.855 2.47 15.855 2.94 19.005 2.94 19.005 2.005 16.385 2.005 16.385 1.315 16.615 1.315 16.615 1.775 19.235 1.775 19.235 3.17 16.515 3.17 16.515 3.75 16.285 3.75 16.285 3.17 15.625 3.17 15.625 2.7 8.45 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 2.215 2.515 2.215 2.515 2.95 5.845 2.95 5.845 2.215 6.075 2.215 6.075 3.27 2.285 3.27  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.27 5.195 2.27 5.195 2.65 2.95 2.65  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 0.845 0.575 0.845 0.575 4.36 0.15 4.36  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.55 1.21 8.945 1.21 8.945 0.845 9.175 0.845 9.175 4.36 8.845 4.36 8.845 1.59 8.55 1.59  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.55 1.595 3.55 1.595 4.59 3.645 4.59 3.645 3.96 3.875 3.96 3.875 4.59 4.385 4.59 4.385 3.96 4.615 3.96 4.615 4.59 7.645 4.59 7.645 3.55 7.875 3.55 7.875 4.59 8.495 4.59 9.52 4.59 9.52 5.49 8.495 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 7.875 0.45 7.875 1.355 7.645 1.355 7.645 0.45 1.595 0.45 1.595 1.35 1.365 1.35 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.285 0.68 6.755 0.68 6.755 1.355 6.525 1.355 6.525 0.91 4.515 0.91 4.515 1.355 4.285 1.355  ;
        POLYGON 2.055 3.5 6.725 3.5 6.725 2.27 7.35 2.27 7.35 2.5 6.955 2.5 6.955 3.73 2.855 3.73 2.855 4.36 2.625 4.36 2.625 3.73 1.825 3.73 1.825 2.555 0.925 2.555 0.925 2.215 1.825 2.215 1.825 1.07 3.85 1.07 3.85 1.3 2.055 1.3  ;
        POLYGON 6.57 3.96 7.185 3.96 7.185 3.09 7.58 3.09 7.58 1.985 5.405 1.985 5.405 1.14 5.635 1.14 5.635 1.755 7.81 1.755 7.81 2.215 8.495 2.215 8.495 2.555 7.81 2.555 7.81 3.32 7.415 3.32 7.415 4.19 6.57 4.19  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.03 2.27 3.84 2.27 3.84 2.94 5.75 2.94 5.75 2.27 7.16 2.27 7.16 2.5 6.01 2.5 6.01 3.17 3.61 3.17 3.61 2.5 3.03 2.5  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 2.15 4.33 2.15 4.33 2.71 4.07 2.71  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 0.77 1.615 0.77 1.615 4.355 1.27 4.355  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.985 0.77 10.49 0.77 10.49 1.59 10.215 1.59 10.215 4.355 9.985 4.355  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.315 4.59 0.315 3.875 0.545 3.875 0.545 4.59 2.455 4.59 2.455 3.875 2.685 3.875 2.685 4.59 4.545 4.59 4.545 3.875 4.775 3.875 4.775 4.59 5.365 4.59 5.365 3.875 5.595 3.875 5.595 4.59 8.865 4.59 8.865 3.875 9.095 3.875 9.095 4.59 9.635 4.59 11.055 4.59 11.055 3.875 11.285 3.875 11.285 4.59 11.76 4.59 11.76 5.49 9.635 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 11.335 0.45 11.335 1.58 11.105 1.58 11.105 0.45 9.095 0.45 9.095 1.58 8.865 1.58 8.865 0.45 2.735 0.45 2.735 1.58 2.505 1.58 2.505 0.45 0.495 0.45 0.495 1.58 0.265 1.58 0.265 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 5.265 0.68 7.735 0.68 7.735 1.11 7.505 1.11 7.505 0.91 5.495 0.91 5.495 1.58 5.265 1.58  ;
        POLYGON 2.015 1.855 2.245 1.855 2.245 2.385 2.8 2.385 2.8 3.4 7.945 3.4 7.945 2.04 4.545 2.04 4.545 0.77 4.775 0.77 4.775 1.81 8.175 1.81 8.175 3.63 3.755 3.63 3.755 4.325 3.525 4.325 3.525 3.63 2.57 3.63 2.57 2.665 2.015 2.665  ;
        POLYGON 7.505 3.875 8.405 3.875 8.405 1.57 6.385 1.57 6.385 1.14 6.615 1.14 6.615 1.34 8.635 1.34 8.635 2.27 9.4 2.27 9.4 1.835 9.635 1.835 9.635 2.645 8.635 2.645 8.635 4.215 7.505 4.215  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.3 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.1 2.215 1.33 2.215 1.33 2.63 3.93 2.63 3.93 2.285 6.45 2.285 6.45 2.63 7.85 2.63 7.85 2.27 9.86 2.27 9.86 2.5 8.08 2.5 8.08 2.86 1.1 2.86  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.3 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 1.825 6.91 1.825 6.91 2.17 7.62 2.17 7.62 2.4 6.68 2.4 6.68 2.055 3.05 2.055 3.05 2.4 1.77 2.4  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5505 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.47 1.365 15.15 1.365 15.15 1.595 12.805 1.595 12.805 2.985 15.1 2.985 15.1 3.215 12.47 3.215  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.6603 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.95 2.96 18.59 2.96 19.075 2.96 19.075 1.79 16.95 1.79 16.95 0.695 17.335 0.695 17.335 1.43 19.345 1.43 19.345 0.695 19.575 0.695 19.575 1.79 19.435 1.79 19.435 4.36 19.205 4.36 19.205 3.32 18.59 3.32 17.235 3.32 17.235 4.36 16.95 4.36  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 2.335 4.59 2.335 3.55 2.565 3.55 2.565 4.59 4.425 4.59 4.425 3.55 4.655 3.55 4.655 4.59 7.915 4.59 7.915 4.01 8.145 4.01 8.145 4.59 11.275 4.59 11.275 4.01 11.505 4.01 11.505 4.59 13.695 4.59 13.695 4.01 13.925 4.01 13.925 4.59 15.885 4.59 15.885 3.55 16.115 3.55 16.115 4.59 18.125 4.59 18.125 3.55 18.355 3.55 18.355 4.59 18.59 4.59 20.335 4.59 20.335 3.55 20.565 3.55 20.565 4.59 21.28 4.59 21.28 5.49 18.59 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.695 0.45 20.695 1.2 20.465 1.2 20.465 0.45 18.455 0.45 18.455 1.2 18.225 1.2 18.225 0.45 16.215 0.45 16.215 1.2 15.985 1.2 15.985 0.675 11.735 0.675 11.735 1.125 11.505 1.125 11.505 0.45 4.655 0.45 4.655 1.595 4.425 1.595 4.425 0.45 0.475 0.45 0.475 1.2 0.245 1.2 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 5.67 0.845 10.49 0.845 10.49 1.075 5.67 1.075  ;
        POLYGON 0.87 3.09 10.09 3.09 10.09 2.27 12.23 2.27 12.23 2.5 10.32 2.5 10.32 3.32 3.635 3.32 3.635 4.36 3.405 4.36 3.405 3.32 1.545 3.32 1.545 4.36 1.315 4.36 1.315 3.32 0.64 3.32 0.64 1.365 2.385 1.365 2.385 0.695 2.615 0.695 2.615 1.595 0.87 1.595  ;
        POLYGON 5.725 3.55 15.38 3.55 15.38 1.135 12.195 1.135 12.195 1.585 6.79 1.585 6.79 1.355 11.965 1.355 11.965 0.905 15.61 0.905 15.61 2.215 18.59 2.215 18.59 2.555 15.61 2.555 15.61 3.78 10.385 3.78 10.385 4.36 10.155 4.36 10.155 3.78 5.955 3.78 5.955 4.36 5.725 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.806 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.15 0.97 2.15 0.97 2.96 0.71 2.96 0.71 2.71 0.115 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.806 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.15 2.715 2.15 2.715 2.71 2.06 2.71 2.06 2.96 1.83 2.96  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 0.845 3.855 0.845 3.855 3.685 3.51 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 4.345 0.475 4.345 0.475 4.59 2.285 4.59 2.285 4.345 2.515 4.345 2.515 4.59 3.175 4.59 4.48 4.59 4.48 5.49 3.175 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 2.735 0.45 2.735 1.165 2.505 1.165 2.505 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.21 3.885 2.945 3.885 2.945 1.625 0.19 1.625 0.19 1.37 0.53 1.37 0.53 1.395 3.175 1.395 3.175 4.115 1.55 4.115 1.55 4.17 1.21 4.17  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.612 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.33 0.71 2.33 0.71 1.905 0.97 1.905 0.97 2.715 0.15 2.715  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.612 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.33 1.83 2.33 1.83 1.9 2.09 1.9 2.09 2.71 1.27 2.71  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.42 0.845 3.77 0.845 3.77 3.685 3.42 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.26 4.59 0.26 3.685 0.49 3.685 0.49 4.59 2.52 4.59 2.52 3.875 2.75 3.875 2.75 4.59 2.97 4.59 4.56 4.59 4.56 3.875 4.79 3.875 4.79 4.59 5.04 4.59 5.04 5.49 2.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 4.77 0.45 4.77 1.165 4.54 1.165 4.54 0.45 2.53 0.45 2.53 1.165 2.3 1.165 2.3 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.28 2.94 2.74 2.94 2.74 1.655 0.26 1.655 0.26 0.845 0.49 0.845 0.49 1.425 2.97 1.425 2.97 3.17 1.51 3.17 1.51 3.75 1.28 3.75  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.205 1.21 2.09 1.21 2.09 2.06 1.205 2.06  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.355 1.77 0.97 1.77 0.97 2.29 4.03 2.29 4.03 2.715 0.355 2.715  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.445 2.79 6.465 2.79 7.485 2.79 7.485 1.6 5.39 1.6 5.39 0.9 8.085 0.9 8.085 3.685 6.465 3.685 5.445 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.875 0.475 3.875 0.475 4.59 2.285 4.59 2.285 3.875 2.515 3.875 2.515 4.59 4.325 4.59 4.325 3.875 4.555 3.875 4.555 4.59 6.465 4.59 6.545 4.59 6.545 4.23 6.775 4.23 6.775 4.59 8.585 4.59 8.585 4.225 8.815 4.225 8.815 4.59 9.52 4.59 9.52 5.49 6.465 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 9.035 0.45 9.035 1.165 8.805 1.165 8.805 0.45 6.85 0.45 6.85 0.64 6.51 0.64 6.51 0.45 4.555 0.45 4.555 1.165 4.325 1.165 4.325 0.45 0.475 0.45 0.475 1.165 0.245 1.165 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.95 4.765 2.95 4.765 1.655 2.32 1.655 2.32 0.845 2.55 0.845 2.55 1.425 4.995 1.425 4.995 1.975 6.465 1.975 6.465 2.315 4.995 2.315 4.995 3.18 3.535 3.18 3.535 3.875 3.305 3.875 3.305 3.18 1.495 3.18 1.495 3.875 1.265 3.875  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.125 2.74 1.145 2.74 1.145 3.345 0.125 3.345  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.82 2.74 2.725 2.74 2.725 3.375 1.82 3.375  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 1.77 2.955 1.77 2.955 2.15 0.565 2.15  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 0.845 4.995 0.845 4.995 3.83 4.63 3.83  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 4.345 1.495 4.345 1.495 4.59 3.645 4.59 3.645 4.345 3.875 4.345 3.875 4.59 4.315 4.59 5.6 4.59 5.6 5.49 4.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 3.875 0.45 3.875 1.35 3.645 1.35 3.645 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.885 3.185 3.885 3.185 0.98 0.475 0.98 0.475 1.355 0.245 1.355 0.245 0.75 3.415 0.75 3.415 1.775 4.315 1.775 4.315 2.115 3.415 2.115 3.415 4.315 2.285 4.315 2.285 4.115 0.475 4.115 0.475 4.315 0.245 4.315  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.16 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.15 0.97 2.15 0.97 2.71 0.115 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 2.15 2.09 2.15 2.09 2.71 1.21 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 2.29 3.21 2.29 3.21 2.71 2.39 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.48 0.845 4.89 0.845 4.89 3.685 4.48 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.32 4.59 1.32 3.875 1.55 3.875 1.55 4.59 3.36 4.59 3.36 3.875 3.59 3.875 3.59 4.59 4.21 4.59 5.58 4.59 5.58 3.875 5.81 3.875 5.81 4.59 6.16 4.59 6.16 5.49 4.21 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.16 -0.45 6.16 0.45 5.83 0.45 5.83 1.165 5.6 1.165 5.6 0.45 3.59 0.45 3.59 1.165 3.36 1.165 3.36 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.3 3.98 3.3 3.98 1.92 0.3 1.92 0.3 0.845 0.53 0.845 0.53 1.69 4.21 1.69 4.21 3.53 2.57 3.53 2.57 4.11 2.34 4.11 2.34 3.53 0.245 3.53  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.2 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.245 1.73 3.115 1.73 3.115 2.15 1.245 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 2.38 3.995 2.38 3.995 1.77 5 1.77 5 2.61 1.79 2.61  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.33 0.995 2.33 0.995 2.84 5.785 2.84 5.785 2.415 6.02 2.415 6.02 3.07 0.15 3.07  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.55 2.925 9.26 2.925 9.58 2.925 9.58 1.6 7.25 1.6 7.25 0.895 9.93 0.895 9.93 3.63 9.26 3.63 7.55 3.63  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.505 0.475 3.505 0.475 4.59 2.285 4.59 2.285 3.975 2.515 3.975 2.515 4.59 4.325 4.59 4.325 3.975 4.555 3.975 4.555 4.59 6.585 4.59 6.585 3.875 6.815 3.875 6.815 4.59 8.625 4.59 8.625 3.875 8.855 3.875 8.855 4.59 9.26 4.59 10.665 4.59 10.665 3.875 10.895 3.875 10.895 4.59 11.2 4.59 11.2 5.49 9.26 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.2 -0.45 11.2 0.45 10.895 0.45 10.895 1.165 10.665 1.165 10.665 0.45 8.71 0.45 8.71 0.64 8.37 0.64 8.37 0.45 6.415 0.45 6.415 1.165 6.185 1.165 6.185 0.45 0.555 0.45 0.555 0.695 0.325 0.695 0.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 3.3 6.625 3.3 6.625 1.625 5.5 1.625 5.5 1.52 3.305 1.52 3.305 0.71 3.535 0.71 3.535 1.29 5.755 1.29 5.755 1.395 6.855 1.395 6.855 1.97 9.26 1.97 9.26 2.31 6.855 2.31 6.855 3.53 5.575 3.53 5.575 4.11 5.345 4.11 5.345 3.53 3.535 3.53 3.535 4.11 3.305 4.11 3.305 3.53 1.495 3.53 1.495 4.11 1.265 4.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.16 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.165 0.975 2.165 0.975 2.71 0.115 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 1.21 2.09 1.21 2.09 2.115 1.23 2.115  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.32 1.21 3.21 1.21 3.21 2.115 2.32 2.115  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.83 2.33 4.5 2.33 4.5 2.71 3.83 2.71  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 2.89 5.235 2.89 5.585 2.89 5.585 0.845 6.045 0.845 6.045 3.685 5.235 3.685 5.19 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.305 4.59 0.305 3.155 0.535 3.155 0.535 4.59 2.345 4.59 2.345 3.155 2.575 3.155 2.575 4.59 4.565 4.59 4.565 4.345 4.795 4.345 4.795 4.59 5.235 4.59 6.16 4.59 6.16 5.49 5.235 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.16 -0.45 6.16 0.45 4.795 0.45 4.795 1.35 4.565 1.35 4.565 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.325 2.695 3.595 2.695 3.595 2.985 4.73 2.985 4.73 2.005 3.44 2.005 3.44 0.98 0.535 0.98 0.535 1.355 0.305 1.355 0.305 0.75 3.67 0.75 3.67 1.775 5.235 1.775 5.235 2.115 4.96 2.115 4.96 3.215 3.365 3.215 3.365 2.925 1.555 2.925 1.555 3.215 1.325 3.215  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.15 0.97 2.15 0.97 2.71 0.115 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 2.15 2.09 2.15 2.09 2.71 1.2 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.32 2.29 3.21 2.29 3.21 2.71 2.32 2.71  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.44 2.33 4.33 2.33 4.33 2.71 3.44 2.71  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 0.845 6.1 0.845 6.1 3.685 5.58 3.685 5.58 1.725 5.19 1.725  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.3 4.59 0.3 3.875 0.53 3.875 0.53 4.59 2.34 4.59 2.34 4.345 2.57 4.345 2.57 4.59 4.38 4.59 4.38 3.875 4.61 3.875 4.61 4.59 5.23 4.59 6.6 4.59 6.6 3.875 6.83 3.875 6.83 4.59 7.28 4.59 7.28 5.49 5.23 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 6.85 0.45 6.85 1.165 6.62 1.165 6.62 0.45 4.61 0.45 4.61 0.695 4.38 0.695 4.38 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.32 3.415 4.56 3.415 4.56 1.6 0.245 1.6 0.245 1.37 4.79 1.37 4.79 2.38 5.23 2.38 5.23 2.72 4.79 2.72 4.79 3.645 3.59 3.645 3.59 4.235 3.36 4.235 3.36 3.765 1.32 3.765  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 13.44 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.79 1.77 3.89 1.77 3.89 2.15 2.79 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.825 2.38 4.52 2.38 4.52 1.77 6.03 1.77 6.03 2.15 4.75 2.15 4.75 2.61 2.825 2.61  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.975 1.21 2.09 1.21 2.09 1.31 6.49 1.31 6.49 1.83 7.105 1.83 7.105 2.06 6.26 2.06 6.26 1.54 2.145 1.54 2.145 2.06 0.975 2.06  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.33 0.97 2.33 0.97 2.84 4.98 2.84 4.98 2.47 8.125 2.47 8.125 2.7 5.21 2.7 5.21 3.07 0.115 3.07  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.54 2.92 10.55 2.92 11.77 2.92 11.77 1.6 9.485 1.6 9.485 0.9 12.21 0.9 12.21 3.64 10.55 3.64 9.54 3.64  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.26 4.59 0.26 3.325 0.49 3.325 0.49 4.59 2.3 4.59 2.3 3.795 2.53 3.795 2.53 4.59 4.34 4.59 4.34 3.795 4.57 3.795 4.57 4.59 6.38 4.59 6.38 3.795 6.61 3.795 6.61 4.59 8.42 4.59 8.42 3.795 8.65 3.795 8.65 4.59 10.55 4.59 10.64 4.59 10.64 3.875 10.87 3.875 10.87 4.59 12.68 4.59 12.68 3.875 12.91 3.875 12.91 4.59 13.44 4.59 13.44 5.49 10.55 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 13.44 -0.45 13.44 0.45 13.13 0.45 13.13 1.165 12.9 1.165 12.9 0.45 10.945 0.45 10.945 0.64 10.605 0.64 10.605 0.45 8.65 0.45 8.65 0.695 8.42 0.695 8.42 0.45 0.49 0.45 0.49 1.165 0.26 1.165 0.26 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.28 3.3 5.4 3.3 5.4 3.2 8.86 3.2 8.86 1.26 6.715 1.26 6.715 1.08 4.285 1.08 4.285 0.85 6.94 0.85 6.94 1.03 9.09 1.03 9.09 1.975 10.55 1.975 10.55 2.315 9.09 2.315 9.09 3.43 7.63 3.43 7.63 4.01 7.4 4.01 7.4 3.43 5.59 3.43 5.59 4.11 5.36 4.11 5.36 3.53 3.55 3.53 3.55 4.11 3.32 4.11 3.32 3.53 1.51 3.53 1.51 4.11 1.28 4.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__antenna
  CLASS core gf180mcu_fd_sc_mcu9t5v0__antennaCELL ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__antenna 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 1.12 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    gf180mcu_fd_sc_mcu9t5v0__antennaDIFFAREA 0.4068 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.315 0.475 1.315 0.475 3.215 0.15 3.215  ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.12 4.59 1.12 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 1.12 -0.45 1.12 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__antenna
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.415 2.655 2.415 2.655 3.27 1.83 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.285 0.97 2.285 0.97 2.71 0.115 2.71  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.805 3.78 1.805 3.78 2.815 2.95 2.815  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 1.77 2.285 1.77 2.285 0.845 2.515 0.845 2.515 2.15 1.495 2.15 1.495 3.685 1.265 3.685  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.515 4.59 3.485 4.59 3.485 3.875 3.715 3.875 3.715 4.59 4.48 4.59 4.48 5.49 2.515 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 3.815 0.45 3.815 1.565 3.585 1.565 3.585 0.45 0.475 0.45 0.475 1.165 0.245 1.165 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.55 0.475 3.55 0.475 4.13 2.285 4.13 2.285 3.55 2.515 3.55 2.515 4.36 0.245 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.755 5.12 1.755 5.12 2.3 4 2.3  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.77 3.66 1.77 3.66 2.56 5.69 2.56 5.69 2.155 6.605 2.155 6.605 2.79 3.41 2.79  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 1.665 0.98 1.665 0.98 2.15 0.115 2.15  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.2876 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.715 3.02 5.86 3.02 5.86 3.83 5.63 3.83 5.63 3.25 3.7 3.25 3.7 3.83 3.45 3.83 3.45 3.25 2.33 3.25 2.33 1.155 1.375 1.155 1.375 0.925 3.01 0.925 3.01 0.68 4.92 0.68 4.92 1.49 2.715 1.49  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.33 4.59 1.33 4.345 1.56 4.345 1.56 4.59 6.88 4.59 7.28 4.59 7.28 5.49 6.88 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 6.88 0.45 6.88 1.165 6.65 1.165 6.65 0.45 2.78 0.45 2.78 0.695 2.55 0.695 2.55 0.45 0.54 0.45 0.54 1.165 0.31 1.165 0.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.31 3.48 2.68 3.48 2.68 4.06 4.61 4.06 4.61 3.48 4.84 3.48 4.84 4.06 6.65 4.06 6.65 3.48 6.88 3.48 6.88 4.29 2.445 4.29 2.445 3.765 0.54 3.765 0.54 4.36 0.31 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 13.44 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.325 5.895 1.325 5.895 2.11 5.665 2.11 5.665 1.57 0.97 1.57 0.97 2.615 1.905 2.615 1.905 2.42 2.135 2.42 2.135 2.845 0.71 2.845  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.96 4.365 1.96 4.365 2.475 8.31 2.475 8.31 2.71 3.43 2.71 3.43 2.19 1.43 2.19 1.43 2.385 1.2 2.385  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.63 2.33 12.47 2.33 12.47 2.15 12.73 2.15 12.73 2.33 12.735 2.33 12.735 2.75 9.63 2.75  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.136 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.41 3.075 7.58 3.075 7.58 3.015 8.55 3.015 8.55 2 6.345 2 6.345 1.095 2.37 1.095 2.37 0.865 6.575 0.865 6.575 1.77 9.605 1.77 9.605 0.84 9.835 0.84 9.835 1.79 11.845 1.79 11.845 0.84 12.075 0.84 12.075 2.02 8.83 2.02 8.83 3.245 7.815 3.245 7.815 3.885 7.585 3.885 7.585 3.305 5.775 3.305 5.775 3.885 5.545 3.885 5.545 3.305 3.735 3.305 3.735 3.835 3.505 3.835 3.505 3.305 1.695 3.305 1.695 3.835 1.41 3.835  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 9.85 4.59 9.85 3.935 10.19 3.935 10.19 4.59 11.89 4.59 11.89 3.935 12.23 3.935 12.23 4.59 13.25 4.59 13.44 4.59 13.44 5.49 13.25 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 13.44 -0.45 13.44 0.45 13.195 0.45 13.195 1.56 12.965 1.56 12.965 0.45 10.955 0.45 10.955 1.56 10.725 1.56 10.725 0.45 8.535 0.45 8.535 1.085 8.305 1.085 8.305 0.45 4.67 0.45 4.67 0.635 4.33 0.635 4.33 0.45 0.695 0.45 0.695 0.69 0.465 0.69 0.465 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.445 3.535 0.675 3.535 0.675 4.115 2.485 4.115 2.485 3.535 2.715 3.535 2.715 4.115 4.525 4.115 4.525 3.535 4.755 3.535 4.755 4.115 6.565 4.115 6.565 3.535 6.795 3.535 6.795 4.115 8.55 4.115 8.55 3.475 13.25 3.475 13.25 4.23 12.91 4.23 12.91 3.705 11.21 3.705 11.21 4.23 10.87 4.23 10.87 3.705 8.88 3.705 8.88 4.345 0.445 4.345  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.93 1.21 3.83 1.21 3.83 2.115 2.93 2.115  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.95 2.33 4.915 2.33 4.915 2.71 3.95 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.25 1.21 2.09 1.21 2.09 2.115 1.25 2.115  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.13 2.175 0.98 2.175 0.98 2.71 0.13 2.71  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 0.845 2.58 0.845 2.58 2.855 3.6 2.855 3.6 3.83 3.365 3.83 3.365 3.355 2.35 3.355  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.33 4.59 1.33 3.875 1.56 3.875 1.56 4.59 4.62 4.59 5.04 4.59 5.04 5.49 4.62 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 4.62 0.45 4.62 1.165 4.39 1.165 4.39 0.45 0.54 0.45 0.54 1.165 0.31 1.165 0.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.31 3.41 2.05 3.41 2.05 4.06 4.39 4.06 4.39 3.48 4.62 3.48 4.62 4.29 1.82 4.29 1.82 3.645 0.54 3.645 0.54 4.36 0.31 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 1.72 7.21 1.72 7.21 2.315 5.75 2.315  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.95 1.83 5.51 1.83 5.51 2.56 7.86 2.56 7.86 2.18 8.27 2.18 8.27 2.79 4.95 2.79  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.22 1.21 2.09 1.21 2.09 2.06 1.65 2.06 1.65 1.63 1.22 1.63  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.69 1.77 0.97 1.77 0.97 2.29 4.03 2.29 4.03 2.52 0.69 2.52  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.3222 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.72 3.02 7.615 3.02 7.615 3.83 7.385 3.83 7.385 3.25 5.575 3.25 5.575 3.83 4.345 3.83 4.345 1.49 4.34 1.49 4.34 1.105 2.55 1.105 2.55 1.49 2.32 1.49 2.32 0.68 2.55 0.68 2.55 0.875 6.365 0.875 6.365 0.68 6.595 0.68 6.595 1.49 6.365 1.49 6.365 1.105 4.72 1.105  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.875 1.495 3.875 1.495 4.59 3.305 4.59 3.305 3.875 3.535 3.875 3.535 4.59 8.635 4.59 8.96 4.59 8.96 5.49 8.635 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 8.635 0.45 8.635 1.165 8.405 1.165 8.405 0.45 4.61 0.45 4.61 0.64 4.27 0.64 4.27 0.45 0.475 0.45 0.475 1.165 0.245 1.165 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.415 4.025 3.415 4.025 4.06 6.365 4.06 6.365 3.48 6.595 3.48 6.595 4.06 8.405 4.06 8.405 3.48 8.635 3.48 8.635 4.29 3.795 4.29 3.795 3.645 2.515 3.645 2.515 4.225 2.285 4.225 2.285 3.645 0.475 3.645 0.475 4.225 0.245 4.225  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.21 2.27 11.66 2.27 11.66 2.63 14.185 2.63 14.185 2.215 14.415 2.215 14.415 2.86 11.44 2.86 11.44 2.71 11.21 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.325 1.77 13.185 1.77 13.185 0.68 16.355 0.68 16.355 2.555 16.125 2.555 16.125 0.91 13.415 0.91 13.415 2.4 12.47 2.4 12.47 2 9.555 2 9.555 2.555 9.325 2.555  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.81 2.27 3.21 2.27 3.21 2.785 4.205 2.785 4.205 2.27 6.07 2.27 6.07 2.5 4.435 2.5 4.435 3.015 2.81 3.015  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 7.715 1.77 7.715 2.215 7.955 2.215 7.955 2.555 7.485 2.555 7.485 2 3.975 2 3.975 2.555 3.745 2.555 3.745 2 0.915 2 0.915 2.555 0.15 2.555  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.095 3.08 11.245 3.08 11.245 3.09 14.765 3.09 14.765 1.14 14.995 1.14 14.995 3.09 16.015 3.09 16.015 3.9 15.27 3.9 15.27 3.32 13.975 3.32 13.975 3.9 13.745 3.9 13.745 3.32 11.935 3.32 11.935 3.9 11.705 3.9 11.705 3.32 11.195 3.32 11.195 3.315 10.965 3.315 10.965 3.31 9.895 3.31 9.895 3.9 8.865 3.9 8.865 1.985 7.945 1.985 7.945 1.54 2.285 1.54 2.285 0.73 2.515 0.73 2.515 1.31 6.365 1.31 6.365 0.73 6.595 0.73 6.595 1.31 8.175 1.31 8.175 1.755 8.865 1.755 8.865 0.73 10.915 0.73 10.915 1.54 9.095 1.54  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.245 1.495 3.245 1.495 4.59 3.305 4.59 3.305 3.705 3.535 3.705 3.535 4.59 5.345 4.59 5.345 3.705 5.575 3.705 5.575 4.59 7.385 4.59 7.385 3.705 7.615 3.705 7.615 4.59 17.035 4.59 17.36 4.59 17.36 5.49 17.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 17.035 0.45 17.035 1.54 16.805 1.54 16.805 0.45 12.955 0.45 12.955 1.54 12.725 1.54 12.725 0.45 8.635 0.45 8.635 1.525 8.405 1.525 8.405 0.45 4.555 0.45 4.555 1.07 4.325 1.07 4.325 0.45 0.475 0.45 0.475 1.54 0.245 1.54 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.785 2.38 2.785 2.38 3.245 8.635 3.245 8.635 4.13 10.685 4.13 10.685 3.54 10.915 3.54 10.915 4.13 12.725 4.13 12.725 3.55 12.955 3.55 12.955 4.13 14.765 4.13 14.765 3.55 14.995 3.55 14.995 4.13 16.805 4.13 16.805 3.245 17.035 3.245 17.035 4.36 8.405 4.36 8.405 3.475 6.595 3.475 6.595 4.055 6.365 4.055 6.365 3.475 4.555 3.475 4.555 4.055 4.325 4.055 4.325 3.475 2.515 3.475 2.515 4.055 2.15 4.055 2.15 3.015 0.475 3.015 0.475 4.055 0.245 4.055  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 1.21 2.695 1.21 2.695 2.115 1.77 2.115  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 1.705 0.97 1.705 0.97 2.595 0.115 2.595  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.925 1.615 3.815 1.615 3.815 2.15 2.925 2.15  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.045 1.615 4.915 1.615 4.915 2.15 4.045 2.15  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 0.75 3.28 0.75 3.28 1.06 4.63 1.06 4.63 0.92 4.86 0.92 4.86 1.29 3.05 1.29 3.05 0.98 1.53 0.98 1.53 3.83 1.27 3.83  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.52 4.59 4.53 4.59 4.53 3.875 4.76 3.875 4.76 4.59 5.6 4.59 5.6 5.49 2.52 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 3.74 0.45 3.74 0.83 3.51 0.83 3.51 0.45 0.48 0.45 0.48 1.3 0.25 1.3 0.25 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 3.55 0.48 3.55 0.48 4.13 2.29 4.13 2.29 3.55 2.52 3.55 2.52 4.36 0.25 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 1.77 2.955 1.77 2.955 2.215 1.765 2.215  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.305 1.155 2.305 1.155 2.445 3.51 2.445 3.51 1.77 3.77 1.77 3.77 2.775 0.63 2.775  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.56 1.725 5.45 1.725 5.45 2.47 8.43 2.47 8.43 2.7 4.56 2.7  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 1.77 7.295 1.77 7.295 2.15 5.75 2.15  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.341 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 3.4 4.07 3.4 4.07 1.525 2.205 1.525 2.205 0.715 2.435 0.715 2.435 1.265 4.73 1.265 4.73 0.93 5.465 0.93 5.465 0.695 5.695 0.695 5.695 0.93 7.705 0.93 7.705 0.79 7.935 0.79 7.935 1.16 4.96 1.16 4.96 1.495 4.33 1.495 4.33 3.63 1.21 3.63  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 6.505 4.59 6.505 4.345 6.735 4.345 6.735 4.59 8.815 4.59 9.52 4.59 9.52 5.49 8.815 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 9.055 0.45 9.055 0.7 8.825 0.7 8.825 0.45 6.815 0.45 6.815 0.7 6.585 0.7 6.585 0.45 4.395 0.45 4.395 0.7 4.165 0.7 4.165 0.45 0.475 0.45 0.475 1.17 0.245 1.17 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.28 0.475 3.28 0.475 3.86 8.585 3.86 8.585 3.28 8.815 3.28 8.815 4.09 0.245 4.09  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.16 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.755 5.805 1.755 5.805 2.17 6.64 2.17 6.64 2.4 5.575 2.4 5.575 1.985 4.89 1.985 4.89 2.15 3.85 2.15 3.85 2.4 3.51 2.4  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.545 2.215 1.775 2.215 1.775 2.63 5.115 2.63 5.115 2.215 5.345 2.215 5.345 2.63 6.87 2.63 6.87 2.215 8.725 2.215 8.725 2.86 1.545 2.86  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.86 2.27 10.2 2.27 10.2 2.73 13.505 2.73 13.505 2.215 13.735 2.215 13.735 2.73 18.96 2.73 18.96 2.27 19.45 2.27 19.45 2.96 9.86 2.96  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.52 1.755 14.42 1.755 14.42 2.27 16.5 2.27 16.5 2.5 14.19 2.5 14.19 2.15 13.96 2.15 13.96 1.985 12.86 1.985 12.86 2.5 12.52 2.5  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.682 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.085 1.31 2.955 1.31 2.955 0.68 3.185 0.68 3.185 1.18 18.67 1.18 18.67 1.525 3.04 1.525 3.04 1.54 1.315 1.54 1.315 3.09 8.285 3.09 8.285 3.9 8.055 3.9 8.055 3.32 6.245 3.32 6.245 3.9 5.75 3.9 5.75 3.32 4.205 3.32 4.205 3.9 3.975 3.9 3.975 3.32 2.165 3.32 2.165 3.9 1.935 3.9 1.935 3.32 1.085 3.32  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 11.475 4.59 11.475 3.65 11.705 3.65 11.705 4.59 16.795 4.59 16.795 3.65 17.025 3.65 17.025 4.59 19.685 4.59 20.16 4.59 20.16 5.49 19.685 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.16 -0.45 20.16 0.45 19.735 0.45 19.735 1.035 19.505 1.035 19.505 0.45 17.34 0.45 17.34 0.95 17 0.95 17 0.45 14.68 0.45 14.68 0.95 14.34 0.95 14.34 0.45 12.02 0.45 12.02 0.95 11.68 0.95 11.68 0.45 9.36 0.45 9.36 0.95 9.02 0.95 9.02 0.45 5.225 0.45 5.225 0.695 4.995 0.695 4.995 0.45 0.905 0.45 0.905 1.165 0.675 1.165 0.675 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.915 3.55 1.145 3.55 1.145 4.13 2.955 4.13 2.955 3.55 3.185 3.55 3.185 4.13 4.995 4.13 4.995 3.55 5.225 3.55 5.225 4.13 7.035 4.13 7.035 3.55 7.265 3.55 7.265 4.13 9.075 4.13 9.075 3.19 19.685 3.19 19.685 4.36 19.455 4.36 19.455 3.42 14.365 3.42 14.365 4.36 14.135 4.36 14.135 3.42 9.305 3.42 9.305 4.36 0.915 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.16 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.145 2.415 5.375 2.415 5.375 2.865 6.04 2.865 6.04 3.27 5.145 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 2.165 4.33 2.165 4.33 2.71 3.45 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.255 1.21 2.09 1.21 2.09 2.065 1.255 2.065  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.135 2.255 1.015 2.255 1.015 2.71 0.135 2.71  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.36 1.67 3.21 1.67 3.21 2.23 2.36 2.23  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.184 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.425 1.075 2.655 1.075 2.655 1.21 5.685 1.21 5.685 0.68 5.915 0.68 5.915 1.59 4.795 1.59 4.795 3.685 4.565 3.685 4.565 1.44 2.425 1.44  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.875 1.595 3.875 1.595 4.59 2.615 4.59 5.815 4.59 6.16 4.59 6.16 5.49 5.815 5.49 2.615 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.16 -0.45 6.16 0.45 3.955 0.45 3.955 0.98 3.725 0.98 3.725 0.45 0.515 0.45 0.515 1.3 0.285 1.3 0.285 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 2.385 2.94 2.385 2.875 2.615 2.875 2.615 3.685 2.385 3.685 2.385 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 3.545 3.55 3.775 3.55 3.775 4.13 5.585 4.13 5.585 3.55 5.815 3.55 5.815 4.36 3.545 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.225 2.47 10.165 2.47 10.165 1.21 10.49 1.21 10.49 2.7 7.225 2.7  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.3 1.21 8.47 1.21 8.47 2.115 8.24 2.115 8.24 1.59 7.3 1.59  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 1.665 3.845 1.665 3.845 2.18 2.945 2.18  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.89 2.44 4.49 2.44 4.49 2.205 5.48 2.205 5.48 2.67 1.89 2.67  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.715 1.915 2.485 1.915 2.485 1.205 4.89 1.205 4.89 1.52 6.37 1.52 6.37 1.75 4.63 1.75 4.63 1.435 2.715 1.435 2.715 2.145 1.01 2.145 1.01 2.785 0.715 2.785  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.11125 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 1.315 0.475 1.315 0.475 1.455 2.025 1.455 2.025 0.745 5.35 0.745 5.35 1.06 6.765 1.06 6.765 0.92 6.995 0.92 6.995 3.02 10.88 3.02 10.88 0.845 11.11 0.845 11.11 3.83 9.76 3.83 9.76 3.25 7.95 3.25 7.95 3.83 7.72 3.83 7.72 3.25 6.765 3.25 6.765 1.29 5.12 1.29 5.12 0.975 2.255 0.975 2.255 1.685 0.245 1.685  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.33 4.59 2.33 4.4 2.67 4.4 2.67 4.59 4.39 4.59 4.39 4.4 4.73 4.4 4.73 4.59 11.065 4.59 11.76 4.59 11.76 5.49 11.065 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 9.15 0.45 9.15 1.3 8.92 1.3 8.92 0.45 5.81 0.45 5.81 0.83 5.58 0.83 5.58 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.9 1.595 2.9 1.595 3.48 3.405 3.48 3.405 2.9 3.635 2.9 3.635 3.48 5.465 3.48 5.465 2.9 5.695 2.9 5.695 3.71 1.365 3.71  ;
        POLYGON 0.345 3.36 0.575 3.36 0.575 3.94 6.665 3.94 6.665 3.48 6.895 3.48 6.895 4.06 8.74 4.06 8.74 3.48 8.97 3.48 8.97 4.06 11.065 4.06 11.065 4.29 6.665 4.29 6.665 4.17 0.345 4.17  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 22.4 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.21 1.91 16.95 1.91 16.95 1.21 18.23 1.21 18.23 1.72 19.77 1.72 19.77 2.37 21.45 2.37 21.45 2.6 19.54 2.6 19.54 1.95 18 1.95 18 1.44 17.27 1.44 17.27 2.4 16.93 2.4 16.93 2.14 14.55 2.14 14.55 2.5 14.21 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.15 2.37 16.7 2.37 16.7 2.63 17.51 2.63 17.51 1.77 17.77 1.77 17.77 2.27 19.31 2.27 19.31 2.5 17.74 2.5 17.74 2.86 16.47 2.86 16.47 2.6 16.15 2.6  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.7 1.855 3.51 1.855 3.51 1.21 3.77 1.21 3.77 1.755 6.425 1.755 6.425 2.37 8.16 2.37 8.16 2.6 6.195 2.6 6.195 1.985 3.925 1.985 3.925 2.4 3.695 2.4 3.695 2.085 1.04 2.085 1.04 2.6 0.7 2.6  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.315 1.985 2.315 1.985 2.63 5.735 2.63 5.735 2.215 5.965 2.215 5.965 2.86 1.27 2.86  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.11 2.27 9.65 2.27 9.65 2.71 9.11 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.0645 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.395 3.05 1.395 3.05 0.735 4.66 0.735 4.66 1.25 8.555 1.25 8.555 0.68 8.785 0.68 8.785 1.25 11.165 1.25 11.165 0.68 11.395 0.68 11.395 1.25 13.405 1.25 13.405 0.68 13.635 0.68 13.635 1.25 16.49 1.25 16.49 0.735 18.69 0.735 18.69 1.26 21.745 1.26 21.745 0.68 21.975 0.68 21.975 1.49 18.46 1.49 18.46 0.965 16.72 0.965 16.72 1.48 13.85 1.48 13.85 3.09 20.955 3.09 20.955 3.9 20.725 3.9 20.725 3.32 18.915 3.32 18.915 3.9 18.685 3.9 18.685 3.32 16.875 3.32 16.875 3.9 16.645 3.9 16.645 3.32 14.835 3.32 14.835 3.9 14.605 3.9 14.605 3.32 13.59 3.32 13.59 1.48 4.43 1.48 4.43 0.965 3.28 0.965 3.28 1.625 0.245 1.625  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.09 0.525 3.09 0.525 4.59 2.335 4.59 2.335 3.55 2.565 3.55 2.565 4.59 4.375 4.59 4.375 3.55 4.605 3.55 4.605 4.59 6.415 4.59 6.415 3.55 6.645 3.55 6.645 4.59 8.455 4.59 8.455 3.55 8.685 3.55 8.685 4.59 21.975 4.59 22.4 4.59 22.4 5.49 21.975 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 22.4 -0.45 22.4 0.45 19.935 0.45 19.935 1.02 19.705 1.02 19.705 0.45 15.855 0.45 15.855 1.02 15.625 1.02 15.625 0.45 12.515 0.45 12.515 1.02 12.285 1.02 12.285 0.45 10.275 0.45 10.275 1.02 10.045 1.02 10.045 0.45 6.645 0.45 6.645 1.02 6.415 1.02 6.415 0.45 2.565 0.45 2.565 1.165 2.335 1.165 2.335 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.315 3.09 10.34 3.09 10.34 3.075 12.465 3.075 12.465 3.9 12.235 3.9 12.235 3.305 10.425 3.305 10.425 3.9 10.195 3.9 10.195 3.32 7.665 3.32 7.665 3.9 7.435 3.9 7.435 3.32 5.625 3.32 5.625 3.9 5.395 3.9 5.395 3.32 3.585 3.32 3.585 3.9 3.355 3.9 3.355 3.32 1.545 3.32 1.545 3.9 1.315 3.9  ;
        POLYGON 9.175 3.55 9.405 3.55 9.405 4.13 11.215 4.13 11.215 3.535 11.445 3.535 11.445 4.13 13.305 4.13 13.305 3.545 13.535 3.545 13.535 4.13 15.625 4.13 15.625 3.55 15.855 3.55 15.855 4.13 17.665 4.13 17.665 3.55 17.895 3.55 17.895 4.13 19.705 4.13 19.705 3.55 19.935 3.55 19.935 4.13 21.745 4.13 21.745 3.09 21.975 3.09 21.975 4.36 9.175 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 2.415 7.725 2.415 7.725 3.27 6.8 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.145 1.77 6.01 1.77 6.01 2.15 5.145 2.15  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.67 1.77 3.83 1.77 3.83 2.15 2.67 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.05 2.255 4.91 2.255 4.91 2.71 4.05 2.71  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.22 1.21 2.145 1.21 2.145 2.06 1.22 2.06  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.235 1.07 2.235 1.07 2.71 0.115 2.71  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.1692 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.22 2.875 6.24 2.875 6.24 1.49 3.16 1.49 3.16 0.68 3.39 0.68 3.39 1.21 7.24 1.21 7.24 0.68 7.47 0.68 7.47 1.59 6.47 1.59 6.47 3.215 6.22 3.215  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.4 4.59 0.4 3.875 0.63 3.875 0.63 4.59 2.44 4.59 2.44 3.875 2.67 3.875 2.67 4.59 7.47 4.59 7.84 4.59 7.84 5.49 7.47 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 5.43 0.45 5.43 0.695 5.2 0.695 5.2 0.45 0.71 0.45 0.71 1.165 0.48 1.165 0.48 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.94 4.465 2.94 4.465 3.81 4.125 3.81 4.125 3.17 1.71 3.17 1.71 3.7 1.365 3.7  ;
        POLYGON 3.16 3.55 3.39 3.55 3.39 4.13 5.2 4.13 5.2 3.55 7.47 3.55 7.47 4.36 3.16 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.7 2.345 11.775 2.345 11.775 1.21 12.96 1.21 12.96 2.575 9.7 2.575  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.945 1.21 11.05 1.21 11.05 2.115 9.945 2.115  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.605 2.38 7.605 2.38 7.605 1.77 8.81 1.77 8.81 2.61 5.605 2.61  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.255 1.77 6.77 1.77 6.77 2.15 5.255 2.15  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.415 4.065 2.415 4.065 2.645 0.97 2.645 0.97 3.27 0.115 3.27  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.77 2.09 1.77 2.09 2.15 0.825 2.15  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.2758 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 0.68 0.51 0.68 0.51 0.925 4.98 0.925 4.98 0.68 5.21 0.68 5.21 0.925 9.16 0.925 9.16 0.845 9.47 0.845 9.47 2.875 13.255 2.875 13.255 0.845 13.485 0.845 13.485 3.105 12.465 3.105 12.465 3.685 12.235 3.685 12.235 3.105 10.425 3.105 10.425 3.685 10.195 3.685 10.195 3.105 9.04 3.105 9.04 1.49 0.28 1.49 0.28 1.01 0.28 0.925  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.28 4.59 0.28 3.875 0.51 3.875 0.51 4.59 2.32 4.59 2.32 3.875 2.55 3.875 2.55 4.59 4.36 4.59 4.36 3.875 4.59 3.875 4.59 4.59 13.485 4.59 14 4.59 14 5.49 13.485 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14 -0.45 14 0.45 11.445 0.45 11.445 0.695 11.215 0.695 11.215 0.45 7.35 0.45 7.35 0.695 7.12 0.695 7.12 0.45 2.55 0.45 2.55 0.695 2.32 0.695 2.32 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.3 2.875 8.37 2.875 8.37 3.685 8.14 3.685 8.14 3.105 6.33 3.105 6.33 3.685 6.1 3.685 6.1 3.105 3.57 3.105 3.57 3.685 3.34 3.685 3.34 3.105 1.53 3.105 1.53 3.685 1.3 3.685  ;
        POLYGON 5.08 3.335 5.31 3.335 5.31 3.915 7.12 3.915 7.12 3.335 7.35 3.335 7.35 3.915 9.16 3.915 9.16 3.335 9.39 3.335 9.39 3.915 11.215 3.915 11.215 3.335 11.445 3.335 11.445 3.915 13.255 3.915 13.255 3.335 13.485 3.335 13.485 4.145 5.08 4.145  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 26.32 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.865 1.755 25.095 1.755 25.095 2.555 24.865 2.555 24.865 1.985 21.015 1.985 21.015 2.4 20.785 2.4 20.785 1.985 19.45 1.985 19.45 2.15 18.095 2.15 18.095 2.555 17.865 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.75 2.27 20.32 2.27 20.32 2.63 22.595 2.63 22.595 2.215 23.055 2.215 23.055 2.77 22.78 2.77 22.78 2.86 20.135 2.86 20.135 2.77 19.75 2.77  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.67 1.37 12.775 1.37 12.775 1.425 16.835 1.425 16.835 2.555 16.605 2.555 16.605 1.655 12.855 1.655 12.855 2.4 12.625 2.4 12.625 1.6 9.93 1.6 9.93 2.555 9.67 2.555  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.69 1.83 12.33 1.83 12.33 2.63 13.955 2.63 13.955 2.54 14.665 2.54 14.665 2.215 14.895 2.215 14.895 2.77 14.14 2.77 14.14 2.86 12.1 2.86 12.1 2.5 11.69 2.5  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.755 8.055 1.755 8.055 2.555 7.825 2.555 7.825 2.15 6.31 2.15 6.31 1.985 3.975 1.985 3.975 2.555 3.745 2.555 3.745 1.985 1.055 1.985 1.055 2.555 0.825 2.555  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.215 3.515 2.215 3.515 2.785 5.49 2.785 5.49 2.625 5.785 2.625 5.785 2.215 6.015 2.215 6.015 2.855 5.71 2.855 5.71 3.015 3.285 3.015 3.285 2.445 2.09 2.445 2.09 2.71 1.83 2.71  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.2844 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 0.91 13.49 0.91 13.49 0.925 24.73 0.925 24.73 0.71 25.73 0.71 25.73 1.195 17.515 1.195 17.515 2.785 17.895 2.785 17.895 3 19.925 3 19.925 3.09 23.035 3.09 23.035 3 24.655 3 24.655 3.9 24.425 3.9 24.425 3.23 23.22 3.23 23.22 3.32 22.615 3.32 22.615 3.9 22.385 3.9 22.385 3.32 20.575 3.32 20.575 3.9 20.345 3.9 20.345 3.32 19.74 3.32 19.74 3.23 18.535 3.23 18.535 3.9 18.305 3.9 18.305 3.23 17.665 3.23 17.665 3.015 17.285 3.015 17.285 1.155 13.405 1.155 13.405 1.14 8.69 1.14 8.69 1.195 0.19 1.195  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.245 0.475 3.245 0.475 4.59 2.285 4.59 2.285 3.705 2.515 3.705 2.515 4.59 4.325 4.59 4.325 3.705 4.555 3.705 4.555 4.59 6.365 4.59 6.365 3.56 6.595 3.56 6.595 4.59 8.405 4.59 8.405 3.545 8.635 3.545 8.635 4.59 25.675 4.59 26.32 4.59 26.32 5.49 25.675 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 26.32 -0.45 26.32 0.45 23.635 0.45 23.635 0.695 23.405 0.695 23.405 0.45 19.555 0.45 19.555 0.695 19.325 0.695 19.325 0.45 15.475 0.45 15.475 0.695 15.245 0.695 15.245 0.45 11.45 0.45 11.45 0.68 11.11 0.68 11.11 0.45 6.65 0.45 6.65 0.68 6.31 0.68 6.31 0.45 2.57 0.45 2.57 0.68 2.23 0.68 2.23 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 3.245 5.93 3.245 5.93 3.085 9.455 3.085 9.455 3.09 14.325 3.09 14.325 3 16.495 3 16.495 3.9 16.265 3.9 16.265 3.23 14.51 3.23 14.51 3.9 14.225 3.9 14.225 3.32 12.415 3.32 12.415 3.9 12.185 3.9 12.185 3.32 10.375 3.32 10.375 3.9 10.145 3.9 10.145 3.32 9.405 3.32 9.405 3.315 7.615 3.315 7.615 4.055 7.385 4.055 7.385 3.315 6.15 3.315 6.15 3.475 5.575 3.475 5.575 4.055 5.345 4.055 5.345 3.475 3.535 3.475 3.535 4.055 3.305 4.055 3.305 3.475 1.495 3.475 1.495 4.055 1.265 4.055  ;
        POLYGON 9.125 3.545 9.355 3.545 9.355 4.13 11.165 4.13 11.165 3.55 11.395 3.55 11.395 4.13 13.205 4.13 13.205 3.55 13.435 3.55 13.435 4.13 15.245 4.13 15.245 3.46 15.475 3.46 15.475 4.13 17.285 4.13 17.285 3.405 17.515 3.405 17.515 4.13 19.325 4.13 19.325 3.46 19.555 3.46 19.555 4.13 21.365 4.13 21.365 3.55 21.595 3.55 21.595 4.13 23.405 4.13 23.405 3.46 23.635 3.46 23.635 4.13 25.445 4.13 25.445 3.245 25.675 3.245 25.675 4.36 9.125 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 3.36 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.015 1.77 1.015 2.71 0.71 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 2.89 2.665 2.89 2.665 1.59 2.39 1.59 2.39 0.74 2.895 0.74 2.895 3.775 2.39 3.775  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.4 1.595 3.4 1.595 4.59 2.215 4.59 3.36 4.59 3.36 5.49 2.215 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 3.36 -0.45 3.36 0.45 1.595 0.45 1.595 1.08 1.365 1.08 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.93 2.94 1.93 1.54 0.245 1.54 0.245 0.74 0.475 0.74 0.475 1.31 2.16 1.31 2.16 1.775 2.215 1.775 2.215 2.585 2.16 2.585 2.16 3.17 0.575 3.17 0.575 3.775 0.345 3.775  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.33 0.63 2.33 0.63 2 0.97 2 0.97 2.71 0.15 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.485 2.73 2.75 2.73 2.98 2.73 2.98 1.59 2.33 1.59 2.33 0.71 2.715 0.71 2.715 1.21 3.28 1.21 3.28 3.015 2.75 3.015 2.715 3.015 2.715 4.36 2.485 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.55 1.495 3.55 1.495 4.59 2.75 4.59 3.505 4.59 3.505 3.55 3.735 3.55 3.735 4.59 4.48 4.59 4.48 5.49 2.75 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 3.835 0.45 3.835 1.52 3.605 1.52 3.605 0.45 1.595 0.45 1.595 1.165 1.365 1.165 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.09 1.2 3.09 1.2 1.625 0.245 1.625 0.245 0.71 0.475 0.71 0.475 1.395 1.43 1.395 1.43 2.27 2.75 2.27 2.75 2.5 1.43 2.5 1.43 3.32 0.475 3.32 0.475 4.36 0.245 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.915 1.77 0.915 2.585 0.41 2.585 0.41 2.71 0.15 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.207 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.675 2.875 3.22 2.875 3.51 2.875 3.51 2 2.675 2 2.675 0.73 2.905 0.73 2.905 1.77 4.915 1.77 4.915 0.73 5.145 0.73 5.145 2 4.005 2 4.005 2.875 5.045 2.875 5.045 3.685 4.815 3.685 4.815 3.105 3.22 3.105 2.905 3.105 2.905 4.36 2.675 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.55 1.495 3.55 1.495 4.59 3.22 4.59 3.695 4.59 3.695 3.55 3.925 3.55 3.925 4.59 5.6 4.59 5.6 5.49 3.22 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.025 0.45 4.025 1.54 3.795 1.54 3.795 0.45 1.785 0.45 1.785 1.165 1.555 1.165 1.555 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.09 1.145 3.09 1.145 1.54 0.245 1.54 0.245 0.73 0.475 0.73 0.475 1.31 1.375 1.31 1.375 2.27 3.22 2.27 3.22 2.5 1.375 2.5 1.375 3.32 0.475 3.32 0.475 4.36 0.245 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_3
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 1.91 2.27 1.91 2.65 0.63 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.605 3.09 4.62 3.09 5.575 3.09 5.575 1.95 3.605 1.95 3.605 0.68 3.865 0.68 3.865 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 4.36 5.745 4.36 5.745 3.32 4.62 3.32 3.835 3.32 3.835 4.36 3.605 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.62 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 7.84 4.59 7.84 5.49 4.62 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 3.09 2.14 3.09 2.14 1.92 1.365 1.92 1.365 0.68 1.595 0.68 1.595 1.69 2.37 1.69 2.37 2.27 4.62 2.27 4.62 2.5 2.37 2.5 2.37 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.215 4.205 2.215 4.205 2.65 0.685 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.845 2.88 8.74 2.88 8.97 2.88 8.97 2.04 5.845 2.04 5.845 0.68 6.075 0.68 6.075 1.72 8.055 1.72 8.055 0.68 8.315 0.68 8.315 1.72 10.325 1.72 10.325 0.68 10.555 0.68 10.555 1.72 12.565 1.72 12.565 0.68 12.795 0.68 12.795 1.985 9.47 1.985 9.47 2.88 12.695 2.88 12.695 4.36 12.465 4.36 12.465 3.32 10.455 3.32 10.455 4.36 10.225 4.36 10.225 3.32 8.74 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 6.075 3.32 6.075 4.36 5.845 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 8.74 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.22 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 14.56 4.59 14.56 5.49 13.22 5.49 8.74 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.165 9.205 1.165 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.975 4.435 2.975 4.435 1.985 1.365 1.985 1.365 0.68 1.595 0.68 1.595 1.755 3.605 1.755 3.605 0.68 3.835 0.68 3.835 1.755 4.665 1.755 4.665 2.27 8.74 2.27 8.74 2.65 4.665 2.65 4.665 3.205 3.735 3.205 3.735 4.36 3.505 4.36 3.505 3.205 1.595 3.205 1.595 4.36 1.365 4.36  ;
        POLYGON 9.7 2.215 13.22 2.215 13.22 2.65 9.7 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_8
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.242 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.13 2.27 5.64 2.27 5.64 2.65 0.13 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.926 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.135 2.84 12.91 2.84 13.5 2.84 13.5 2.04 8.135 2.04 8.135 0.68 8.365 0.68 8.365 1.755 10.375 1.755 10.375 0.68 10.605 0.68 10.605 1.755 12.385 1.755 12.385 0.68 12.845 0.68 12.845 1.755 14.855 1.755 14.855 0.68 15.085 0.68 15.085 1.755 17.095 1.755 17.095 0.68 17.325 0.68 17.325 1.755 19.335 1.755 19.335 0.68 19.565 0.68 19.565 1.985 14 1.985 14 2.84 19.465 2.84 19.465 4.36 19.235 4.36 19.235 3.32 17.225 3.32 17.225 4.36 16.995 4.36 16.995 3.32 14.985 3.32 14.985 4.36 14.755 4.36 14.755 3.32 12.91 3.32 12.745 3.32 12.745 4.36 12.515 4.36 12.515 3.32 10.505 3.32 10.505 4.36 10.275 4.36 10.275 3.32 8.365 3.32 8.365 4.36 8.135 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 2.435 4.59 2.435 3.55 2.665 3.55 2.665 4.59 4.675 4.59 4.675 3.55 4.905 3.55 4.905 4.59 6.915 4.59 6.915 3.55 7.145 3.55 7.145 4.59 9.155 4.59 9.155 3.875 9.385 3.875 9.385 4.59 11.395 4.59 11.395 3.55 11.625 3.55 11.625 4.59 12.91 4.59 13.635 4.59 13.635 3.55 13.865 3.55 13.865 4.59 15.875 4.59 15.875 3.55 16.105 3.55 16.105 4.59 18.115 4.59 18.115 3.55 18.345 3.55 18.345 4.59 19.63 4.59 20.355 4.59 20.355 3.55 20.585 3.55 20.585 4.59 21.28 4.59 21.28 5.49 19.63 5.49 12.91 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.685 0.45 20.685 1.49 20.455 1.49 20.455 0.45 18.445 0.45 18.445 1.49 18.215 1.49 18.215 0.45 16.205 0.45 16.205 1.49 15.975 1.49 15.975 0.45 13.965 0.45 13.965 1.49 13.735 1.49 13.735 0.45 11.725 0.45 11.725 1.49 11.495 1.49 11.495 0.45 9.485 0.45 9.485 1.49 9.255 1.49 9.255 0.45 7.245 0.45 7.245 1.49 7.015 1.49 7.015 0.45 5.005 0.45 5.005 1.49 4.775 1.49 4.775 0.45 2.765 0.45 2.765 1.49 2.535 1.49 2.535 0.45 0.525 0.45 0.525 1.49 0.295 1.49 0.295 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.415 2.88 5.895 2.88 5.895 2.04 1.415 2.04 1.415 0.68 1.645 0.68 1.645 1.72 3.655 1.72 3.655 0.68 3.885 0.68 3.885 1.72 5.895 1.72 5.895 0.68 6.225 0.68 6.225 2.27 12.91 2.27 12.91 2.5 6.225 2.5 6.225 4.36 5.82 4.36 5.82 3.32 3.785 3.32 3.785 4.36 3.555 4.36 3.555 3.32 1.645 3.32 1.645 4.36 1.415 4.36  ;
        POLYGON 14.23 2.215 19.63 2.215 19.63 2.555 14.23 2.555  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_12
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.656 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.44 2.27 7.83 2.27 7.83 2.65 0.44 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.568 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.325 2.96 16.98 2.96 17.805 2.96 17.805 2.04 10.325 2.04 10.325 0.68 10.555 0.68 10.555 1.72 12.565 1.72 12.565 0.68 12.795 0.68 12.795 1.72 14.805 1.72 14.805 0.68 15.035 0.68 15.035 1.72 17.045 1.72 17.045 0.68 17.305 0.68 17.305 1.72 19.285 1.72 19.285 0.68 19.515 0.68 19.515 1.72 21.525 1.72 21.525 0.68 21.755 0.68 21.755 1.72 23.765 1.72 23.765 0.68 23.995 0.68 23.995 1.72 26.005 1.72 26.005 0.68 26.235 0.68 26.235 1.985 18.555 1.985 18.555 2.96 26.065 2.96 26.135 2.96 26.135 4.36 26.065 4.36 25.905 4.36 25.905 3.32 23.895 3.32 23.895 4.36 23.665 4.36 23.665 3.32 21.655 3.32 21.655 4.36 21.425 4.36 21.425 3.32 19.415 3.32 19.415 4.36 19.185 4.36 19.185 3.32 17.175 3.32 17.175 4.36 16.98 4.36 16.945 4.36 16.945 3.32 14.935 3.32 14.935 4.36 14.705 4.36 14.705 3.32 12.695 3.32 12.695 4.36 12.465 4.36 12.465 3.32 10.555 3.32 10.555 4.36 10.325 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 16.98 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 20.305 4.59 20.305 3.55 20.535 3.55 20.535 4.59 22.545 4.59 22.545 3.55 22.775 3.55 22.775 4.59 24.785 4.59 24.785 3.55 25.015 3.55 25.015 4.59 26.065 4.59 27.025 4.59 27.025 3.55 27.255 3.55 27.255 4.59 28 4.59 28 5.49 26.065 5.49 16.98 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 28 -0.45 28 0.45 27.355 0.45 27.355 1.49 27.125 1.49 27.125 0.45 25.115 0.45 25.115 1.49 24.885 1.49 24.885 0.45 22.875 0.45 22.875 1.49 22.645 1.49 22.645 0.45 20.635 0.45 20.635 1.49 20.405 1.49 20.405 0.45 18.395 0.45 18.395 1.49 18.165 1.49 18.165 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.88 8.06 2.88 8.06 2.04 1.365 2.04 1.365 0.68 1.595 0.68 1.595 1.72 3.605 1.72 3.605 0.68 3.835 0.68 3.835 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 1.72 8.085 1.72 8.085 0.68 8.425 0.68 8.425 2.27 16.98 2.27 16.98 2.63 8.425 2.63 8.425 4.36 8.06 4.36 8.06 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 18.785 2.215 26.065 2.215 26.065 2.555 18.785 2.555  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_16
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 34.72 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.07 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.215 9.845 2.215 9.845 2.65 0.685 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 18.21 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.565 2.885 21.1 2.885 22.285 2.885 22.285 2.03 12.565 2.03 12.565 0.68 12.825 0.68 12.825 1.72 14.805 1.72 14.805 0.68 15.035 0.68 15.035 1.72 17.045 1.72 17.045 0.68 17.275 0.68 17.275 1.72 19.285 1.72 19.285 0.68 19.515 0.68 19.515 1.72 21.525 1.72 21.525 0.68 21.755 0.68 21.755 1.72 23.765 1.72 23.765 0.68 23.995 0.68 23.995 1.72 26.005 1.72 26.005 0.68 26.235 0.68 26.235 1.72 28.245 1.72 28.245 0.68 28.475 0.68 28.475 1.72 30.485 1.72 30.485 0.68 30.715 0.68 30.715 1.72 32.725 1.72 32.725 0.68 32.955 0.68 32.955 1.98 23.035 1.98 23.035 2.88 32.425 2.88 32.855 2.88 32.855 4.36 32.625 4.36 32.625 3.32 32.425 3.32 30.615 3.32 30.615 4.36 30.385 4.36 30.385 3.32 28.375 3.32 28.375 4.36 28.145 4.36 28.145 3.32 26.135 3.32 26.135 4.36 25.905 4.36 25.905 3.32 23.895 3.32 23.895 4.36 23.665 4.36 23.665 3.32 21.655 3.32 21.655 4.36 21.425 4.36 21.425 3.32 21.1 3.32 19.415 3.32 19.415 4.36 19.185 4.36 19.185 3.32 17.175 3.32 17.175 4.36 16.945 4.36 16.945 3.32 14.935 3.32 14.935 4.36 14.705 4.36 14.705 3.32 12.795 3.32 12.795 4.36 12.565 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.875 11.575 3.875 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 20.305 4.59 20.305 3.55 20.535 3.55 20.535 4.59 21.1 4.59 22.545 4.59 22.545 3.55 22.775 3.55 22.775 4.59 24.785 4.59 24.785 3.55 25.015 3.55 25.015 4.59 27.025 4.59 27.025 3.55 27.255 3.55 27.255 4.59 29.265 4.59 29.265 3.55 29.495 3.55 29.495 4.59 31.505 4.59 31.505 3.55 31.735 3.55 31.735 4.59 32.425 4.59 33.745 4.59 33.745 3.55 33.975 3.55 33.975 4.59 34.72 4.59 34.72 5.49 32.425 5.49 21.1 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 34.72 -0.45 34.72 0.45 34.075 0.45 34.075 1.49 33.845 1.49 33.845 0.45 31.835 0.45 31.835 1.49 31.605 1.49 31.605 0.45 29.595 0.45 29.595 1.49 29.365 1.49 29.365 0.45 27.355 0.45 27.355 1.49 27.125 1.49 27.125 0.45 25.115 0.45 25.115 1.49 24.885 1.49 24.885 0.45 22.875 0.45 22.875 1.49 22.645 1.49 22.645 0.45 20.635 0.45 20.635 1.49 20.405 1.49 20.405 0.45 18.395 0.45 18.395 1.49 18.165 1.49 18.165 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.9 10.225 2.9 10.225 1.975 1.365 1.975 1.365 0.68 1.595 0.68 1.595 1.72 3.605 1.72 3.605 0.68 3.835 0.68 3.835 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 1.72 8.085 1.72 8.085 0.68 8.315 0.68 8.315 1.72 10.325 1.72 10.325 0.68 10.555 0.68 10.555 2.27 21.1 2.27 21.1 2.65 10.555 2.65 10.555 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 23.265 2.215 32.425 2.215 32.425 2.65 23.265 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_20
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.698 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.33 2.09 2.33 2.09 2.71 0.87 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.849 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.745 4.99 1.745 4.99 2.15 4.63 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.64 0.84 7.13 0.84 7.13 1.65 6.87 1.65 6.87 3.685 6.64 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.635 1.595 3.635 1.595 4.59 5.44 4.59 5.44 3.875 5.67 3.875 5.67 4.59 6.345 4.59 6.385 4.59 7.28 4.59 7.28 5.49 6.385 5.49 6.345 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 5.89 0.45 5.89 0.69 5.66 0.69 5.66 0.45 1.595 0.45 1.595 1.425 1.365 1.425 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.315 0.475 1.315 0.475 1.83 2.86 1.83 2.86 2.815 2.895 2.815 2.895 3.155 2.63 3.155 2.63 2.06 0.575 2.06 0.575 4.285 0.245 4.285  ;
        POLYGON 2.385 3.475 2.615 3.475 2.615 4.055 4.17 4.055 4.17 1.6 3.55 1.6 3.55 1.37 4.4 1.37 4.4 2.47 6.345 2.47 6.345 2.7 4.65 2.7 4.65 4.285 2.385 4.285  ;
        POLYGON 2.485 0.72 5.43 0.72 5.43 0.92 6.385 0.92 6.385 2.055 5.305 2.055 5.305 1.115 3.32 1.115 3.32 1.83 3.635 1.83 3.635 3.815 3.405 3.815 3.405 2.06 3.09 2.06 3.09 0.95 2.715 0.95 2.715 1.425 2.485 1.425  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.4 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.88 2.33 2.09 2.33 2.09 2.715 0.88 2.715  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.125 2.285 5.465 2.285 5.465 2.71 5.125 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.705 0.84 7.13 0.84 7.13 3.72 6.705 3.72  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.375 4.59 1.375 3.845 1.605 3.845 1.605 4.59 5.685 4.59 5.685 3.88 5.915 3.88 5.915 4.59 6.355 4.59 6.41 4.59 7.725 4.59 7.725 3.88 7.955 3.88 7.955 4.59 8.4 4.59 8.4 5.49 6.41 5.49 6.355 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.4 -0.45 8.4 0.45 8.155 0.45 8.155 1.16 7.925 1.16 7.925 0.45 5.915 0.45 5.915 1.16 5.685 1.16 5.685 0.45 1.605 0.45 1.605 1.165 1.375 1.165 1.375 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.255 0.845 0.485 0.845 0.485 1.83 2.55 1.83 2.55 2.415 3.715 2.415 3.715 2.645 2.32 2.645 2.32 2.06 0.585 2.06 0.585 3.685 0.255 3.685  ;
        POLYGON 2.925 2.875 3.155 2.875 3.155 3.455 4.665 3.455 4.665 1.655 3.615 1.655 3.615 1.315 4.895 1.315 4.895 3.275 6.125 3.275 6.125 2.45 6.355 2.45 6.355 3.505 4.89 3.505 4.89 3.685 2.925 3.685  ;
        POLYGON 2.495 0.68 5.355 0.68 5.355 1.825 6.41 1.825 6.41 2.055 5.125 2.055 5.125 1.085 3.385 1.085 3.385 1.955 4.175 1.955 4.175 3.215 3.945 3.215 3.945 2.185 3.155 2.185 3.155 1.49 2.495 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.64 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.33 2.09 2.33 2.09 2.71 0.87 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.547 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 1.75 6.115 1.75 6.115 2.15 5.75 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9952 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.895 2.91 9.045 2.91 9.045 1.65 7.865 1.65 7.865 0.84 8.095 0.84 8.095 1.39 10.105 1.39 10.105 0.84 10.335 0.84 10.335 1.65 9.39 1.65 9.39 2.91 10.165 2.91 10.165 3.72 9.935 3.72 9.935 3.14 8.125 3.14 8.125 3.72 7.895 3.72  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.845 1.595 3.845 1.595 4.59 4.655 4.59 4.655 4.035 4.885 4.035 4.885 4.59 6.695 4.59 6.695 3.565 6.925 3.565 6.925 4.59 7.665 4.59 8.915 4.59 8.915 3.88 9.145 3.88 9.145 4.59 10.64 4.59 10.64 5.49 7.665 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.64 -0.45 10.64 0.45 9.215 0.45 9.215 1.16 8.985 1.16 8.985 0.45 6.85 0.45 6.85 0.68 6.51 0.68 6.51 0.45 4.61 0.45 4.61 0.68 4.27 0.68 4.27 0.45 1.595 0.45 1.595 1.165 1.365 1.165 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.83 2.55 1.83 2.55 2.47 3.65 2.47 3.65 2.7 2.32 2.7 2.32 2.06 0.575 2.06 0.575 3.685 0.245 3.685  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.91 6.575 0.91 6.575 1.825 7.665 1.825 7.665 2.055 6.345 2.055 6.345 1.14 3.32 1.14 3.32 1.83 4.165 1.83 4.165 3.215 3.935 3.215 3.935 2.06 3.09 2.06 3.09 1.49 2.485 1.49  ;
        POLYGON 2.915 2.93 3.145 2.93 3.145 3.51 5.675 3.51 5.675 2.695 5.29 2.695 5.29 1.6 3.55 1.6 3.55 1.37 5.52 1.37 5.52 2.465 7.665 2.465 7.665 2.695 5.905 2.695 5.905 3.74 2.915 3.74  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_3
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.33 2.09 2.33 2.09 2.71 0.87 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.735 1.77 6.115 1.77 6.115 2.15 5.735 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.2448 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.785 2.97 8.56 2.97 8.96 2.97 8.96 1.62 7.685 1.62 7.685 0.68 7.915 0.68 7.915 1.39 9.925 1.39 9.925 0.68 10.155 0.68 10.155 1.62 9.42 1.62 9.42 2.97 10.055 2.97 10.055 3.78 9.825 3.78 9.825 3.2 8.56 3.2 8.015 3.2 8.015 3.78 7.785 3.78  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.845 1.595 3.845 1.595 4.59 4.725 4.59 4.725 4.35 4.955 4.35 4.955 4.59 6.765 4.59 6.765 3.88 6.995 3.88 6.995 4.59 8.56 4.59 8.805 4.59 8.805 3.88 9.035 3.88 9.035 4.59 10.845 4.59 10.845 3.88 11.075 3.88 11.075 4.59 11.76 4.59 11.76 5.49 8.56 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 11.275 0.45 11.275 1.16 11.045 1.16 11.045 0.45 9.035 0.45 9.035 1.16 8.805 1.16 8.805 0.45 6.85 0.45 6.85 0.635 6.51 0.635 6.51 0.45 4.61 0.45 4.61 0.635 4.27 0.635 4.27 0.45 1.595 0.45 1.595 1.165 1.365 1.165 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.83 2.55 1.83 2.55 2.47 3.65 2.47 3.65 2.7 2.32 2.7 2.32 2.06 0.575 2.06 0.575 3.685 0.245 3.685  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.91 6.575 0.91 6.575 1.85 8.56 1.85 8.56 2.08 6.345 2.08 6.345 1.14 3.32 1.14 3.32 1.83 4.165 1.83 4.165 3.215 3.935 3.215 3.935 2.06 3.09 2.06 3.09 1.49 2.485 1.49  ;
        POLYGON 2.915 2.93 3.145 2.93 3.145 3.51 4.395 3.51 4.395 1.6 3.55 1.6 3.55 1.37 4.625 1.37 4.625 2.505 8.56 2.505 8.56 2.735 5.975 2.735 5.975 3.72 5.745 3.72 5.745 2.735 4.625 2.735 4.625 3.74 2.915 3.74  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 18.48 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.15 1.53 2.15 1.53 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.768 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.175 1.77 8.81 1.77 8.81 2.15 7.175 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.4896 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.015 3.08 14.895 3.08 15.76 3.08 15.76 1.595 10.115 1.595 10.115 0.865 16.835 0.865 16.835 0.84 17.065 0.84 17.065 1.65 16.365 1.65 16.365 3.835 14.895 3.835 10.015 3.835  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.845 1.495 3.845 1.495 4.59 4.915 4.59 4.915 3.88 5.145 3.88 5.145 4.59 6.955 4.59 6.955 3.88 7.185 3.88 7.185 4.59 8.995 4.59 8.995 3.88 9.225 3.88 9.225 4.59 11.035 4.59 11.035 4.35 11.265 4.35 11.265 4.59 13.075 4.59 13.075 4.35 13.305 4.35 13.305 4.59 14.895 4.59 15.115 4.59 15.115 4.35 15.345 4.35 15.345 4.59 17.155 4.59 17.155 3.88 17.385 3.88 17.385 4.59 18.48 4.59 18.48 5.49 14.895 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 18.48 -0.45 18.48 0.45 18.185 0.45 18.185 1.16 17.955 1.16 17.955 0.45 16 0.45 16 0.635 15.66 0.635 15.66 0.45 13.76 0.45 13.76 0.635 13.42 0.635 13.42 0.45 11.52 0.45 11.52 0.635 11.18 0.635 11.18 0.45 9.225 0.45 9.225 0.69 8.995 0.69 8.995 0.45 6.985 0.45 6.985 0.69 6.755 0.69 6.755 0.45 4.61 0.45 4.61 0.625 4.27 0.625 4.27 0.45 1.595 0.45 1.595 0.695 1.365 0.695 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.315 2.035 1.315 2.035 2.47 3.65 2.47 3.65 2.7 1.805 2.7 1.805 1.545 0.475 1.545 0.475 3.685 0.245 3.685  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.855 5.865 0.855 5.865 1.26 7.875 1.26 7.875 0.68 8.105 0.68 8.105 1.26 9.665 1.26 9.665 1.825 14.325 1.825 14.325 2.15 9.435 2.15 9.435 1.49 5.635 1.49 5.635 1.085 3.375 1.085 3.375 2.01 4.175 2.01 4.175 3.685 3.945 3.685 3.945 2.24 3.145 2.24 3.145 1.49 2.485 1.49  ;
        POLYGON 2.925 3.335 3.155 3.335 3.155 3.915 4.405 3.915 4.405 1.78 3.605 1.78 3.605 1.315 3.835 1.315 3.835 1.55 4.635 1.55 4.635 2.91 9.435 2.91 9.435 2.41 14.895 2.41 14.895 2.75 9.665 2.75 9.665 3.14 8.205 3.14 8.205 3.83 7.975 3.83 7.975 3.25 4.635 3.25 4.635 4.145 2.925 4.145  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_8
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 25.2 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.33 1.575 2.33 1.575 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.152 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.04 1.77 11.05 1.77 11.05 2.15 6.04 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.7344 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.255 3.365 21.21 3.365 22.08 3.365 22.08 1.6 12.355 1.6 12.355 0.865 23.785 0.865 23.785 1.65 22.685 1.65 22.685 4.175 21.21 4.175 12.255 4.175  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.505 4.59 1.505 3.845 1.735 3.845 1.735 4.59 5.115 4.59 5.115 3.88 5.345 3.88 5.345 4.59 7.155 4.59 7.155 3.88 7.385 3.88 7.385 4.59 9.195 4.59 9.195 3.88 9.425 3.88 9.425 4.59 11.235 4.59 11.235 3.88 11.465 3.88 11.465 4.59 13.22 4.59 13.22 4.405 13.56 4.405 13.56 4.59 15.26 4.59 15.26 4.405 15.6 4.405 15.6 4.59 17.3 4.59 17.3 4.405 17.64 4.405 17.64 4.59 19.34 4.59 19.34 4.405 19.68 4.405 19.68 4.59 21.21 4.59 21.38 4.59 21.38 4.405 21.72 4.405 21.72 4.59 23.475 4.59 23.475 3.88 23.705 3.88 23.705 4.59 25.2 4.59 25.2 5.49 21.21 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 25.2 -0.45 25.2 0.45 24.905 0.45 24.905 1.16 24.675 1.16 24.675 0.45 22.72 0.45 22.72 0.635 22.38 0.635 22.38 0.45 20.48 0.45 20.48 0.635 20.14 0.635 20.14 0.45 18.24 0.45 18.24 0.635 17.9 0.635 17.9 0.45 16 0.45 16 0.635 15.66 0.635 15.66 0.45 13.76 0.45 13.76 0.635 13.42 0.635 13.42 0.45 11.52 0.45 11.52 0.635 11.18 0.635 11.18 0.45 9.28 0.45 9.28 0.635 8.94 0.635 8.94 0.45 7.04 0.45 7.04 0.635 6.7 0.635 6.7 0.45 4.61 0.45 4.61 0.625 4.27 0.625 4.27 0.45 1.595 0.45 1.595 0.695 1.365 0.695 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.485 2.94 1.805 2.94 1.805 1.6 0.19 1.6 0.19 1.37 2.035 1.37 2.035 2.94 3.365 2.94 3.365 2.415 3.595 2.415 3.595 3.17 0.715 3.17 0.715 3.75 0.485 3.75  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.855 5.865 0.855 5.865 0.865 7.875 0.865 7.875 0.68 8.105 0.68 8.105 1.26 10.115 1.26 10.115 0.68 10.345 0.68 10.345 1.26 11.905 1.26 11.905 1.83 21.035 1.83 21.035 2.15 11.675 2.15 11.675 1.49 5.635 1.49 5.635 1.085 3.375 1.085 3.375 1.955 4.175 1.955 4.175 3.215 3.945 3.215 3.945 2.185 3.145 2.185 3.145 1.49 2.485 1.49  ;
        POLYGON 2.925 3.445 4.405 3.445 4.405 1.655 3.605 1.655 3.605 1.315 4.635 1.315 4.635 2.91 11.465 2.91 11.465 2.45 21.21 2.45 21.21 2.79 11.695 2.79 11.695 3.14 10.445 3.14 10.445 3.94 10.215 3.94 10.215 3.36 4.635 3.36 4.635 3.675 3.155 3.675 3.155 4.255 2.925 4.255  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_12
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 31.92 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 2.33 1.575 2.33 1.575 2.71 0.545 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.536 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.3 2.15 12.125 2.15 12.125 2.71 5.3 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.9792 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.52 3.365 27.62 3.365 27.775 3.365 28.53 3.365 28.53 1.635 14.595 1.635 14.595 0.865 30.505 0.865 30.505 1.65 29.09 1.65 29.09 4.175 27.775 4.175 27.62 4.175 14.52 4.175  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.505 4.59 1.505 3.845 1.735 3.845 1.735 4.59 4.86 4.59 4.86 4.37 5.2 4.37 5.2 4.59 6.9 4.59 6.9 4.37 7.24 4.37 7.24 4.59 8.94 4.59 8.94 4.37 9.28 4.37 9.28 4.59 11.28 4.59 11.28 4.37 11.62 4.37 11.62 4.59 13.5 4.59 13.5 4.405 13.84 4.405 13.84 4.59 15.54 4.59 15.54 4.405 15.88 4.405 15.88 4.59 17.58 4.59 17.58 4.405 17.92 4.405 17.92 4.59 19.62 4.59 19.62 4.405 19.96 4.405 19.96 4.59 21.66 4.59 21.66 4.405 22 4.405 22 4.59 23.7 4.59 23.7 4.405 24.04 4.405 24.04 4.59 25.74 4.59 25.74 4.405 26.08 4.405 26.08 4.59 27.62 4.59 27.775 4.59 27.78 4.59 27.78 4.405 28.12 4.405 28.12 4.59 29.875 4.59 29.875 3.88 30.105 3.88 30.105 4.59 31.92 4.59 31.92 5.49 27.775 5.49 27.62 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 31.92 -0.45 31.92 0.45 31.625 0.45 31.625 1.16 31.395 1.16 31.395 0.45 29.44 0.45 29.44 0.635 29.1 0.635 29.1 0.45 27.2 0.45 27.2 0.635 26.86 0.635 26.86 0.45 24.96 0.45 24.96 0.635 24.62 0.635 24.62 0.45 22.72 0.45 22.72 0.635 22.38 0.635 22.38 0.45 20.48 0.45 20.48 0.635 20.14 0.635 20.14 0.45 18.24 0.45 18.24 0.635 17.9 0.635 17.9 0.45 16 0.45 16 0.635 15.66 0.635 15.66 0.45 13.78 0.45 13.78 0.635 13.405 0.635 13.405 0.45 11.52 0.45 11.52 0.635 11.18 0.635 11.18 0.45 9.28 0.45 9.28 0.635 8.94 0.635 8.94 0.45 7.04 0.45 7.04 0.635 6.7 0.635 6.7 0.45 4.61 0.45 4.61 0.625 4.27 0.625 4.27 0.45 1.595 0.45 1.595 0.695 1.365 0.695 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.485 2.94 1.805 2.94 1.805 1.6 0.19 1.6 0.19 1.37 2.035 1.37 2.035 2.94 3.365 2.94 3.365 2.415 3.595 2.415 3.595 3.17 0.715 3.17 0.715 3.75 0.485 3.75  ;
        POLYGON 2.925 3.445 4.405 3.445 4.405 1.655 3.605 1.655 3.605 1.315 4.635 1.315 4.635 3.33 12.355 3.33 12.355 2.47 27.62 2.47 27.62 2.755 12.7 2.755 12.7 4.14 2.925 4.14  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.855 5.865 0.855 5.865 0.865 14.145 0.865 14.145 1.865 27.775 1.865 27.775 2.16 13.855 2.16 13.855 1.65 5.635 1.65 5.635 1.085 3.375 1.085 3.375 1.955 4.175 1.955 4.175 3.215 3.945 3.215 3.945 2.185 3.145 2.185 3.145 1.49 2.485 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_16
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 3.36 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6765 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.74 1.015 1.74 1.015 2.55 0.71 2.55  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1572 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.21 2.665 1.21 2.665 0.71 2.895 0.71 2.895 3.775 2.565 3.775 2.565 1.59 2.39 1.59  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.24 1.595 3.24 1.595 4.59 2.215 4.59 3.36 4.59 3.36 5.49 2.215 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 3.36 -0.45 3.36 0.45 1.595 0.45 1.595 1.05 1.365 1.05 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.78 1.93 2.78 1.93 1.51 0.245 1.51 0.245 0.71 0.475 0.71 0.475 1.28 2.16 1.28 2.16 1.74 2.215 1.74 2.215 3.01 0.575 3.01 0.575 3.775 0.345 3.775  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.353 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2 0.97 2 0.97 3.27 0.63 3.27  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.5506 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.665 3.96 2.88 3.96 2.88 1.215 2.33 1.215 2.33 0.71 3.11 0.71 3.11 4.3 2.665 4.3  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.96 1.495 3.96 1.495 4.59 2.65 4.59 3.685 4.59 3.685 3.55 3.915 3.55 3.915 4.59 4.48 4.59 4.48 5.49 2.65 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 4.015 0.45 4.015 1.215 3.785 1.215 3.785 0.45 1.595 0.45 1.595 1.215 1.365 1.215 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.5 1.37 3.5 1.37 1.77 0.245 1.77 0.245 0.875 0.475 0.875 0.475 1.54 1.6 1.54 1.6 2.27 2.65 2.27 2.65 2.5 1.6 2.5 1.6 3.73 0.475 3.73 0.475 4.36 0.245 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.035 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.805 1.77 1.53 1.77 1.53 2.215 1.975 2.215 1.975 2.555 0.805 2.555  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.329 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 2.96 4.745 2.96 5.75 2.96 5.75 1.875 3.785 1.875 3.785 1.075 4.015 1.075 4.015 1.645 5.75 1.645 5.75 1.075 6.255 1.075 6.255 4.23 5.925 4.23 5.925 3.19 4.745 3.19 4.015 3.19 4.015 4.23 3.785 4.23  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.42 0.475 3.42 0.475 4.59 2.385 4.59 2.385 3.42 2.615 3.42 2.615 4.59 4.745 4.59 4.805 4.59 4.805 3.42 5.035 3.42 5.035 4.59 7.045 4.59 7.045 3.42 7.275 3.42 7.275 4.59 7.84 4.59 7.84 5.49 4.745 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 7.375 0.45 7.375 1.415 7.145 1.415 7.145 0.45 5.135 0.45 5.135 1.415 4.905 1.415 4.905 0.45 2.895 0.45 2.895 1.415 2.665 1.415 2.665 0.45 0.475 0.45 0.475 1.415 0.245 1.415 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.96 2.205 2.96 2.205 1.36 1.31 1.36 1.31 1.13 2.435 1.13 2.435 2.215 4.745 2.215 4.745 2.555 2.435 2.555 2.435 3.19 1.595 3.19 1.595 4.23 1.365 4.23  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_3
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.706 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.805 1.77 1.53 1.77 1.53 2.215 1.975 2.215 1.975 2.555 0.805 2.555  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.1012 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 3.09 4.745 3.09 5.75 3.09 5.75 1.675 3.785 1.675 3.785 0.875 4.015 0.875 4.015 1.445 5.75 1.445 5.75 0.875 6.255 0.875 6.255 1.875 6.155 1.875 6.155 4.36 5.925 4.36 5.925 3.32 4.745 3.32 4.015 3.32 4.015 4.36 3.785 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.745 4.59 4.805 4.59 4.805 3.55 5.035 3.55 5.035 4.59 7.045 4.59 7.045 3.55 7.275 3.55 7.275 4.59 7.84 4.59 7.84 5.49 4.745 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 7.375 0.45 7.375 1.215 7.145 1.215 7.145 0.45 5.135 0.45 5.135 1.215 4.905 1.215 4.905 0.45 2.895 0.45 2.895 1.215 2.665 1.215 2.665 0.45 0.475 0.45 0.475 1.215 0.245 1.215 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 3.09 2.205 3.09 2.205 1.16 1.31 1.16 1.31 0.93 2.435 0.93 2.435 2.215 4.745 2.215 4.745 2.555 2.435 2.555 2.435 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.412 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 2.215 4.205 2.215 4.205 2.65 0.65 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.2024 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.025 3.09 8.92 3.09 9.15 3.09 9.15 1.745 6.025 1.745 6.025 0.945 6.255 0.945 6.255 1.515 8.265 1.515 8.265 0.945 8.495 0.945 8.495 1.515 10.505 1.515 10.505 0.945 10.735 0.945 10.735 1.515 12.745 1.515 12.745 0.945 12.975 0.945 12.975 1.745 9.65 1.745 9.65 3.09 12.875 3.09 12.875 4.36 12.645 4.36 12.645 3.32 10.635 3.32 10.635 4.36 10.23 4.36 10.23 3.32 8.92 3.32 8.395 3.32 8.395 4.36 8.165 4.36 8.165 3.32 6.255 3.32 6.255 4.36 6.025 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.875 4.855 3.875 4.855 4.59 7.045 4.59 7.045 3.55 7.275 3.55 7.275 4.59 8.92 4.59 9.285 4.59 9.285 3.55 9.515 3.55 9.515 4.59 11.525 4.59 11.525 3.55 11.755 3.55 11.755 4.59 13.51 4.59 13.765 4.59 13.765 3.55 13.995 3.55 13.995 4.59 14.56 4.59 14.56 5.49 13.51 5.49 8.92 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 14.095 0.45 14.095 1.285 13.865 1.285 13.865 0.45 11.855 0.45 11.855 1.215 11.625 1.215 11.625 0.45 9.615 0.45 9.615 1.215 9.385 1.215 9.385 0.45 7.375 0.45 7.375 1.285 7.145 1.285 7.145 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 3.09 4.435 3.09 4.435 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 4.665 1.515 4.665 2.27 8.92 2.27 8.92 2.65 4.665 2.65 4.665 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 9.88 2.27 13.51 2.27 13.51 2.65 9.88 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.118 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.275 1.77 6.01 1.77 6.01 2.215 6.675 2.215 6.675 2.555 1.275 2.555  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.3036 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.485 3.09 13.205 3.09 13.465 3.09 13.465 1.54 8.485 1.54 8.485 1.18 8.715 1.18 8.715 1.31 10.725 1.31 10.725 0.74 10.955 0.74 10.955 1.31 12.965 1.31 12.965 0.74 13.195 0.74 13.195 1.31 15.205 1.31 15.205 0.74 15.435 0.74 15.435 1.31 17.445 1.31 17.445 0.74 17.675 0.74 17.675 1.31 19.685 1.31 19.685 1.18 19.915 1.18 19.915 1.54 14.35 1.54 14.35 3.09 19.815 3.09 19.815 4.36 19.585 4.36 19.585 3.32 17.575 3.32 17.575 4.36 17.345 4.36 17.345 3.32 15.335 3.32 15.335 4.36 14.71 4.36 14.71 3.32 13.205 3.32 13.095 3.32 13.095 4.36 12.865 4.36 12.865 3.32 10.855 3.32 10.855 4.36 10.625 4.36 10.625 3.32 8.715 3.32 8.715 4.36 8.485 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.465 4.59 0.465 3.55 0.695 3.55 0.695 4.59 2.605 4.59 2.605 3.55 2.835 3.55 2.835 4.59 4.845 4.59 4.845 3.55 5.075 3.55 5.075 4.59 7.365 4.59 7.365 3.875 7.595 3.875 7.595 4.59 9.505 4.59 9.505 3.55 9.735 3.55 9.735 4.59 11.745 4.59 11.745 3.55 11.975 3.55 11.975 4.59 13.205 4.59 13.985 4.59 13.985 3.55 14.215 3.55 14.215 4.59 16.225 4.59 16.225 3.55 16.455 3.55 16.455 4.59 18.465 4.59 18.465 3.55 18.695 3.55 18.695 4.59 19.98 4.59 20.705 4.59 20.705 3.55 20.935 3.55 20.935 4.59 21.28 4.59 21.28 5.49 19.98 5.49 13.205 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 21.035 0.45 21.035 1.08 20.805 1.08 20.805 0.45 18.795 0.45 18.795 1.08 18.565 1.08 18.565 0.45 16.555 0.45 16.555 1.08 16.325 1.08 16.325 0.45 14.315 0.45 14.315 1.08 14.085 1.08 14.085 0.45 12.075 0.45 12.075 1.08 11.845 1.08 11.845 0.45 9.835 0.45 9.835 1.08 9.605 1.08 9.605 0.45 7.415 0.45 7.415 1.08 7.185 1.08 7.185 0.45 5.175 0.45 5.175 1.08 4.945 1.08 4.945 0.45 2.935 0.45 2.935 1.08 2.705 1.08 2.705 0.45 0.475 0.45 0.475 1.315 0.245 1.315 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.585 3.09 6.905 3.09 6.905 1.54 1.585 1.54 1.585 1.11 1.815 1.11 1.815 1.31 3.825 1.31 3.825 1.11 4.055 1.11 4.055 1.31 6.065 1.31 6.065 1.11 6.295 1.11 6.295 1.31 7.135 1.31 7.135 2.215 13.205 2.215 13.205 2.555 7.135 2.555 7.135 3.32 6.195 3.32 6.195 4.36 5.965 4.36 5.965 3.32 3.955 3.32 3.955 4.36 3.725 4.36 3.725 3.32 1.815 3.32 1.815 4.36 1.585 4.36  ;
        POLYGON 14.58 2.215 19.98 2.215 19.98 2.555 14.58 2.555  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.824 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.125 7.965 2.125 7.965 2.84 0.685 2.84  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.4048 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.505 3.09 17.105 3.09 17.985 3.09 17.985 1.895 10.505 1.895 10.505 0.945 10.735 0.945 10.735 1.515 12.745 1.515 12.745 0.945 12.975 0.945 12.975 1.665 14.985 1.665 14.985 0.945 15.215 0.945 15.215 1.665 17.225 1.665 17.225 0.945 17.455 0.945 17.455 1.515 19.465 1.515 19.465 0.945 19.695 0.945 19.695 1.515 21.705 1.515 21.705 0.945 21.935 0.945 21.935 1.515 23.945 1.515 23.945 0.945 24.175 0.945 24.175 1.515 26.185 1.515 26.185 0.945 26.415 0.945 26.415 1.745 18.735 1.745 18.735 3.09 26.245 3.09 26.315 3.09 26.315 4.36 26.245 4.36 26.085 4.36 26.085 3.32 24.075 3.32 24.075 4.36 23.845 4.36 23.845 3.32 21.835 3.32 21.835 4.36 21.605 4.36 21.605 3.32 19.595 3.32 19.595 4.36 19.365 4.36 19.365 3.32 17.355 3.32 17.355 4.36 17.125 4.36 17.125 3.32 17.105 3.32 15.115 3.32 15.115 4.36 14.885 4.36 14.885 3.32 12.875 3.32 12.875 4.36 12.645 4.36 12.645 3.32 10.735 3.32 10.735 4.36 10.505 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.875 9.335 3.875 9.335 4.59 11.525 4.59 11.525 3.55 11.755 3.55 11.755 4.59 13.765 4.59 13.765 3.55 13.995 3.55 13.995 4.59 16.005 4.59 16.005 3.55 16.235 3.55 16.235 4.59 17.105 4.59 18.245 4.59 18.245 3.55 18.475 3.55 18.475 4.59 20.485 4.59 20.485 3.55 20.715 3.55 20.715 4.59 22.725 4.59 22.725 3.55 22.955 3.55 22.955 4.59 24.965 4.59 24.965 3.55 25.195 3.55 25.195 4.59 26.245 4.59 27.205 4.59 27.205 3.55 27.435 3.55 27.435 4.59 28 4.59 28 5.49 26.245 5.49 17.105 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 28 -0.45 28 0.45 27.535 0.45 27.535 1.285 27.305 1.285 27.305 0.45 25.295 0.45 25.295 1.215 25.065 1.215 25.065 0.45 23.055 0.45 23.055 1.215 22.825 1.215 22.825 0.45 20.815 0.45 20.815 1.285 20.585 1.285 20.585 0.45 18.575 0.45 18.575 1.215 18.345 1.215 18.345 0.45 16.335 0.45 16.335 1.215 16.105 1.215 16.105 0.45 14.095 0.45 14.095 1.285 13.865 1.285 13.865 0.45 11.855 0.45 11.855 1.285 11.625 1.285 11.625 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 3.09 8.32 3.09 8.32 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.55 0.945 8.55 2.215 17.105 2.215 17.105 2.555 8.55 2.555 8.55 4.36 8.085 4.36 8.085 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 18.965 2.215 26.245 2.215 26.245 2.555 18.965 2.555  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 34.72 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.53 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.215 9.845 2.215 9.845 2.65 0.685 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 15.506 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.745 3.09 21.225 3.09 22.465 3.09 22.465 1.745 12.745 1.745 12.745 0.945 13.005 0.945 13.005 1.515 14.985 1.515 14.985 0.945 15.215 0.945 15.215 1.515 17.225 1.515 17.225 0.945 17.455 0.945 17.455 1.515 19.465 1.515 19.465 0.945 19.695 0.945 19.695 1.515 21.705 1.515 21.705 0.945 21.935 0.945 21.935 1.445 23.945 1.445 23.945 0.945 24.175 0.945 24.175 1.445 26.185 1.445 26.185 0.945 26.415 0.945 26.415 1.445 28.425 1.445 28.425 0.945 28.655 0.945 28.655 1.445 30.665 1.445 30.665 0.945 30.895 0.945 30.895 1.445 32.905 1.445 32.905 0.945 33.135 0.945 33.135 1.675 23.215 1.675 23.215 3.09 32.605 3.09 33.035 3.09 33.035 4.36 32.805 4.36 32.805 3.32 32.605 3.32 30.795 3.32 30.795 4.36 30.565 4.36 30.565 3.32 28.555 3.32 28.555 4.36 28.325 4.36 28.325 3.32 26.315 3.32 26.315 4.36 26.085 4.36 26.085 3.32 24.075 3.32 24.075 4.36 23.845 4.36 23.845 3.32 21.835 3.32 21.835 4.36 21.605 4.36 21.605 3.32 21.225 3.32 19.595 3.32 19.595 4.36 19.365 4.36 19.365 3.32 17.355 3.32 17.355 4.36 17.125 4.36 17.125 3.32 15.115 3.32 15.115 4.36 14.885 4.36 14.885 3.32 12.975 3.32 12.975 4.36 12.745 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.875 11.575 3.875 11.575 4.59 13.765 4.59 13.765 3.55 13.995 3.55 13.995 4.59 16.005 4.59 16.005 3.55 16.235 3.55 16.235 4.59 18.245 4.59 18.245 3.55 18.475 3.55 18.475 4.59 20.485 4.59 20.485 3.55 20.715 3.55 20.715 4.59 21.225 4.59 22.725 4.59 22.725 3.55 22.955 3.55 22.955 4.59 24.965 4.59 24.965 3.55 25.195 3.55 25.195 4.59 27.205 4.59 27.205 3.55 27.435 3.55 27.435 4.59 29.445 4.59 29.445 3.55 29.675 3.55 29.675 4.59 31.685 4.59 31.685 3.55 31.915 3.55 31.915 4.59 32.605 4.59 33.925 4.59 33.925 3.55 34.155 3.55 34.155 4.59 34.72 4.59 34.72 5.49 32.605 5.49 21.225 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 34.72 -0.45 34.72 0.45 34.255 0.45 34.255 1.285 34.025 1.285 34.025 0.45 32.015 0.45 32.015 1.215 31.785 1.215 31.785 0.45 29.775 0.45 29.775 1.215 29.545 1.215 29.545 0.45 27.535 0.45 27.535 1.215 27.305 1.215 27.305 0.45 25.295 0.45 25.295 1.215 25.065 1.215 25.065 0.45 23.055 0.45 23.055 1.215 22.825 1.215 22.825 0.45 20.815 0.45 20.815 1.215 20.585 1.215 20.585 0.45 18.575 0.45 18.575 1.285 18.345 1.285 18.345 0.45 16.335 0.45 16.335 1.285 16.105 1.285 16.105 0.45 14.095 0.45 14.095 1.285 13.865 1.285 13.865 0.45 11.675 0.45 11.675 1.285 11.445 1.285 11.445 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 3.09 10.225 3.09 10.225 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.315 0.945 8.315 1.515 10.325 1.515 10.325 0.945 10.555 0.945 10.555 2.215 21.225 2.215 21.225 2.65 10.455 2.65 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 23.445 2.215 32.605 2.215 32.605 2.65 23.445 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.24 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.353 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.83 0.71 1.83 0.71 1.21 0.97 1.21 0.97 2.53 0.63 2.53  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1264 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 0.945 1.595 0.945 1.595 4.36 1.265 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.24 4.59 2.24 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.24 -0.45 2.24 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 3.36 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.706 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 2.27 1.64 2.27 1.64 2.71 0.36 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.5142 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.55 1.83 3.55 1.83 2.89 1.87 2.89 1.87 2.04 1.365 2.04 1.365 0.945 1.595 0.945 1.595 1.81 2.1 1.81 2.1 3.83 1.595 3.83 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 3.36 4.59 3.36 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 3.36 -0.45 3.36 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.059 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.215 1.83 2.215 1.83 1.77 2.09 1.77 2.09 2.215 2.325 2.215 2.325 2.71 0.685 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.6406 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 3.51 3.09 3.51 1.44 1.365 1.44 1.365 0.68 1.595 0.68 1.595 1.21 3.605 1.21 3.605 0.68 3.835 0.68 3.835 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.48 4.59 4.48 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 2.715 0.45 2.715 0.98 2.485 0.98 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_3
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.412 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 2.38 2.27 2.38 2.65 0.63 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.0284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 2.95 3.09 2.95 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.6 1.515 3.6 0.945 3.835 0.945 3.835 4.36 3.5 4.36 3.5 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 5.6 4.59 5.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.824 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.265 4.26 2.265 4.26 2.645 0.63 2.645  ;
        POLYGON 5.36 2.215 8.88 2.215 8.88 2.65 5.36 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.0568 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 4.63 3.09 4.63 1.745 1.365 1.745 1.365 0.945 1.625 0.945 1.625 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.315 0.945 8.315 1.745 5.13 1.745 5.13 3.09 8.215 3.09 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 10.08 4.59 10.08 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_8
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 16.236 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 6.14 2.27 6.14 2.65 0.63 2.65  ;
        POLYGON 7.66 2.27 13.17 2.27 13.17 2.65 7.66 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.0852 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 6.37 3.09 6.37 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.315 0.945 8.315 1.515 10.325 1.515 10.325 0.945 10.555 0.945 10.555 1.515 12.565 1.515 12.565 0.945 12.795 0.945 12.795 1.745 7.12 1.745 7.12 3.09 12.695 3.09 12.695 4.36 12.465 4.36 12.465 3.32 10.455 3.32 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 14.56 4.59 14.56 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 13.915 0.45 13.915 1.285 13.685 1.285 13.685 0.45 11.675 0.45 11.675 1.285 11.445 1.285 11.445 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_12
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 21.648 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 8.02 2.27 8.02 2.65 0.63 2.65  ;
        POLYGON 9.295 2.27 16.685 2.27 16.685 2.65 9.295 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.1136 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 8.265 3.09 8.265 1.745 1.365 1.745 1.365 0.945 1.625 0.945 1.625 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.315 0.945 8.315 1.515 10.325 1.515 10.325 0.945 10.555 0.945 10.555 1.515 12.565 1.515 12.565 0.945 12.795 0.945 12.795 1.515 14.805 1.515 14.805 0.945 15.035 0.945 15.035 1.515 17.045 1.515 17.045 0.945 17.275 0.945 17.275 1.745 9.065 1.745 9.065 3.09 17.175 3.09 17.175 4.36 16.945 4.36 16.945 3.32 14.935 3.32 14.935 4.36 14.705 4.36 14.705 3.32 12.695 3.32 12.695 4.36 12.465 4.36 12.465 3.32 10.455 3.32 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 19.04 4.59 19.04 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 18.395 0.45 18.395 1.285 18.165 1.285 18.165 0.45 16.155 0.45 16.155 1.285 15.925 1.285 15.925 0.45 13.915 0.45 13.915 1.285 13.685 1.285 13.685 0.45 11.675 0.45 11.675 1.285 11.445 1.285 11.445 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_16
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 27.06 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 9.9 2.27 9.9 2.65 0.63 2.65  ;
        POLYGON 11.11 2.27 20.38 2.27 20.38 2.65 11.11 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 15.142 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 10.13 3.09 10.13 1.745 1.365 1.745 1.365 0.945 1.625 0.945 1.625 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.315 0.945 8.315 1.515 10.325 1.515 10.325 0.945 10.555 0.945 10.555 1.515 12.565 1.515 12.565 0.945 12.795 0.945 12.795 1.515 14.805 1.515 14.805 0.945 15.035 0.945 15.035 1.515 17.045 1.515 17.045 0.945 17.275 0.945 17.275 1.515 19.285 1.515 19.285 0.945 19.515 0.945 19.515 1.515 21.525 1.515 21.525 0.945 21.755 0.945 21.755 1.745 10.88 1.745 10.88 3.09 21.655 3.09 21.655 4.36 21.425 4.36 21.425 3.32 19.415 3.32 19.415 4.36 19.185 4.36 19.185 3.32 17.175 3.32 17.175 4.36 16.945 4.36 16.945 3.32 14.935 3.32 14.935 4.36 14.705 4.36 14.705 3.32 12.695 3.32 12.695 4.36 12.465 4.36 12.465 3.32 10.455 3.32 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 20.305 4.59 20.305 3.55 20.535 3.55 20.535 4.59 22.545 4.59 22.545 3.55 22.775 3.55 22.775 4.59 23.52 4.59 23.52 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 22.875 0.45 22.875 1.285 22.645 1.285 22.645 0.45 20.635 0.45 20.635 1.285 20.405 1.285 20.405 0.45 18.395 0.45 18.395 1.285 18.165 1.285 18.165 0.45 16.155 0.45 16.155 1.285 15.925 1.285 15.925 0.45 13.915 0.45 13.915 1.285 13.685 1.285 13.685 0.45 11.675 0.45 11.675 1.285 11.445 1.285 11.445 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_20
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 16.8 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 2.33 4.33 2.33 4.33 2.71 3.45 2.71  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.57 2.235 1.57 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 1.315 15.055 1.315 15.055 3.215 14.71 3.215  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.61 3.535 3.61 3.535 4.59 6.17 4.59 7.405 4.59 7.405 3.14 7.635 3.14 7.635 4.59 9.195 4.59 12.545 4.59 12.545 3.905 12.775 3.905 12.775 4.59 15.515 4.59 15.845 4.59 15.845 3.875 16.075 3.875 16.075 4.59 16.8 4.59 16.8 5.49 15.515 5.49 9.195 5.49 6.17 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 16.8 -0.45 16.8 0.45 16.175 0.45 16.175 1.165 15.945 1.165 15.945 0.45 12.995 0.45 12.995 0.625 12.765 0.625 12.765 0.45 7.855 0.45 7.855 0.625 7.625 0.625 7.625 0.45 3.435 0.45 3.435 1.13 3.205 1.13 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.425 2.97 4.56 2.97 4.56 1.36 4.325 1.36 4.325 1.02 4.79 1.02 4.79 3.78 4.425 3.78  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 2.99 3.995 2.99 3.995 4.125 6.17 4.125 6.17 4.355 3.765 4.355 3.765 3.22 2.385 3.22  ;
        POLYGON 5.445 1.02 5.675 1.02 5.675 2.05 8.285 2.05 8.285 1.94 8.515 1.94 8.515 2.28 5.675 2.28 5.675 3.78 5.445 3.78  ;
        POLYGON 6.965 2.51 8.965 2.51 8.965 1.315 9.195 1.315 9.195 3.78 8.965 3.78 8.965 2.85 6.965 2.85  ;
        POLYGON 6.125 0.855 9.35 0.855 9.35 0.68 10.775 0.68 10.775 2.3 11.25 2.3 11.25 2.53 10.545 2.53 10.545 1.085 6.355 1.085 6.355 1.82 6.125 1.82  ;
        POLYGON 10.085 1.315 10.315 1.315 10.315 2.76 13.41 2.76 13.41 2.99 10.315 2.99 10.315 3.78 10.085 3.78  ;
        POLYGON 12.05 2.23 14.105 2.23 14.105 1.315 14.48 1.315 14.48 2.455 14.155 2.455 14.155 3.215 13.925 3.215 13.925 2.46 12.05 2.46  ;
        POLYGON 11.47 3.445 15.285 3.445 15.285 1.085 11.655 1.085 11.655 1.225 11.425 1.225 11.425 0.855 15.515 0.855 15.515 3.675 11.47 3.675  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.69 4.325 1.69 4.325 2.235 3.4 2.235  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.33 1.865 2.33 1.865 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.71 1.37 16.09 1.37 16.09 3.27 15.82 3.27 15.82 1.6 15.71 1.6  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.655 4.59 1.655 3.425 1.885 3.425 1.885 4.59 2.325 4.59 3.495 4.59 3.495 3.615 3.725 3.615 3.725 4.59 6.69 4.59 7.925 4.59 7.925 3.145 8.155 3.145 8.155 4.59 9.495 4.59 12.805 4.59 12.805 4.345 13.035 4.345 13.035 4.59 14.8 4.59 14.8 4.345 15.03 4.345 15.03 4.59 16.55 4.59 16.84 4.59 16.84 3.875 17.07 3.875 17.07 4.59 17.36 4.59 17.36 5.49 16.55 5.49 9.495 5.49 6.69 5.49 2.325 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 17.115 0.45 17.115 1.165 16.885 1.165 16.885 0.45 14.93 0.45 14.93 0.64 14.59 0.64 14.59 0.45 13.035 0.45 13.035 1.165 12.805 1.165 12.805 0.45 8.155 0.45 8.155 1.19 7.925 1.19 7.925 0.45 3.625 0.45 3.625 1.19 3.395 1.19 3.395 0.45 1.785 0.45 1.785 1.225 1.555 1.225 1.555 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.635 2.94 2.095 2.94 2.095 1.74 0.435 1.74 0.435 1.315 0.665 1.315 0.665 1.51 2.325 1.51 2.325 3.17 0.865 3.17 0.865 3.75 0.635 3.75  ;
        POLYGON 4.515 2.975 4.56 2.975 4.56 1.08 4.79 1.08 4.79 3.785 4.515 3.785  ;
        POLYGON 2.675 1.315 2.905 1.315 2.905 2.985 4.185 2.985 4.185 4.13 6.69 4.13 6.69 4.36 3.955 4.36 3.955 3.215 2.675 3.215  ;
        POLYGON 5.965 1.08 6.195 1.08 6.195 2.055 8.595 2.055 8.595 2.395 8.365 2.395 8.365 2.285 6.195 2.285 6.195 3.785 5.965 3.785  ;
        POLYGON 7.485 2.515 7.715 2.515 7.715 2.625 8.945 2.625 8.945 2.055 9.265 2.055 9.265 1.315 9.495 1.315 9.495 2.285 9.175 2.285 9.175 3.785 8.945 3.785 8.945 2.855 7.485 2.855  ;
        POLYGON 6.59 1.595 8.805 1.595 8.805 0.68 11.4 0.68 11.4 2.19 11.55 2.19 11.55 2.42 11.17 2.42 11.17 0.91 9.035 0.91 9.035 1.825 6.59 1.825  ;
        POLYGON 10.385 1.315 10.615 1.315 10.615 2.65 13.19 2.65 13.19 2.47 13.53 2.47 13.53 2.88 10.615 2.88 10.615 3.785 10.385 3.785  ;
        POLYGON 12.31 1.92 13.87 1.92 13.87 1.37 14.21 1.37 14.21 1.83 15.525 1.83 15.525 2.06 14.055 2.06 14.055 3.215 13.825 3.215 13.825 2.15 12.31 2.15  ;
        POLYGON 11.785 3.11 12.015 3.11 12.015 3.69 16.32 3.69 16.32 1.14 13.64 1.14 13.64 1.625 11.63 1.625 11.63 1.37 11.97 1.37 11.97 1.395 13.41 1.395 13.41 0.91 16.55 0.91 16.55 3.92 11.785 3.92  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.6 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.43 2.33 4.33 2.33 4.33 2.71 3.43 2.71  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.33 1.705 2.33 1.705 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.71 2.89 17.555 2.89 17.785 2.89 17.785 1.64 15.71 1.64 15.71 1.37 18.29 1.37 18.29 3.23 17.555 3.23 15.71 3.23  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.495 4.59 1.495 3.425 1.725 3.425 1.725 4.59 2.165 4.59 3.435 4.59 3.435 3.515 3.665 3.515 3.665 4.59 6.3 4.59 7.535 4.59 7.535 3.045 7.765 3.045 7.765 4.59 9.265 4.59 12.805 4.59 12.805 4.345 13.035 4.345 13.035 4.59 14.745 4.59 14.745 4.345 14.975 4.345 14.975 4.59 16.785 4.59 16.785 4.345 17.015 4.345 17.015 4.59 18.75 4.59 18.825 4.59 18.825 4.345 19.055 4.345 19.055 4.59 19.6 4.59 19.6 5.49 18.75 5.49 9.265 5.49 6.3 5.49 2.165 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.6 -0.45 19.6 0.45 19.355 0.45 19.355 1.165 19.125 1.165 19.125 0.45 17.17 0.45 17.17 0.64 16.83 0.64 16.83 0.45 14.93 0.45 14.93 0.64 14.59 0.64 14.59 0.45 13.09 0.45 13.09 0.64 12.75 0.64 12.75 0.45 7.985 0.45 7.985 0.625 7.755 0.625 7.755 0.45 3.565 0.45 3.565 1.145 3.335 1.145 3.335 0.45 1.725 0.45 1.725 1.225 1.495 1.225 1.495 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.94 1.935 2.94 1.935 2.005 0.375 2.005 0.375 1.315 0.605 1.315 0.605 1.775 2.165 1.775 2.165 3.17 0.705 3.17 0.705 3.75 0.475 3.75  ;
        POLYGON 4.555 2.875 4.56 2.875 4.56 1.375 4.455 1.375 4.455 1.035 4.79 1.035 4.79 3.685 4.555 3.685  ;
        POLYGON 2.515 1.315 2.845 1.315 2.845 2.985 4.125 2.985 4.125 4.03 6.3 4.03 6.3 4.26 3.895 4.26 3.895 3.215 2.515 3.215  ;
        POLYGON 5.575 1.035 5.805 1.035 5.805 2.01 8.355 2.01 8.355 1.9 8.585 1.9 8.585 2.24 5.805 2.24 5.805 3.685 5.575 3.685  ;
        POLYGON 7.04 2.47 9.035 2.47 9.035 1.315 9.265 1.315 9.265 3.685 9.03 3.685 9.03 2.7 7.04 2.7  ;
        POLYGON 6.2 0.855 9.42 0.855 9.42 0.68 11.395 0.68 11.395 2.755 11.165 2.755 11.165 1.085 6.54 1.085 6.54 1.78 6.2 1.78  ;
        POLYGON 10.155 1.315 10.385 1.315 10.385 2.985 11.625 2.985 11.625 2.47 13.53 2.47 13.53 2.7 11.855 2.7 11.855 3.215 10.385 3.215 10.385 3.685 10.155 3.685  ;
        POLYGON 12.31 1.92 13.87 1.92 13.87 1.37 14.21 1.37 14.21 1.87 17.555 1.87 17.555 2.21 14.055 2.21 14.055 3.215 13.825 3.215 13.825 2.15 12.31 2.15  ;
        POLYGON 11.73 3.5 18.52 3.5 18.52 1.14 11.915 1.14 11.915 1.49 11.685 1.49 11.685 0.68 11.915 0.68 11.915 0.91 18.75 0.91 18.75 3.73 11.73 3.73  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.31 3.77 2.31 3.77 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.03 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.59 1.21 13.91 1.21 13.91 2.025 13.59 2.025  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.665 2.235 1.575 2.235 1.575 2.71 0.665 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.83 3.45 15.93 3.45 16.16 3.45 16.16 0.845 16.39 0.845 16.39 3.83 15.93 3.83 15.83 3.83  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.305 4.59 1.305 3.425 1.535 3.425 1.535 4.59 2.035 4.59 3.045 4.59 3.045 3.515 3.275 3.515 3.275 4.59 5.755 4.59 7.125 4.59 7.125 3.515 7.355 3.515 7.355 4.59 8.375 4.59 8.865 4.59 8.865 3.355 9.095 3.355 9.095 4.59 9.59 4.59 10.115 4.59 13.185 4.59 13.185 4.26 13.525 4.26 13.525 4.59 14.95 4.59 15.28 4.59 15.28 3.735 15.51 3.735 15.51 4.59 15.93 4.59 17.18 4.59 17.18 3.875 17.41 3.875 17.41 4.59 17.92 4.59 17.92 5.49 15.93 5.49 14.95 5.49 10.115 5.49 9.59 5.49 8.375 5.49 5.755 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.51 0.45 17.51 1.165 17.28 1.165 17.28 0.45 13.25 0.45 13.25 1.225 13.02 1.225 13.02 0.45 8.475 0.45 8.475 1.225 8.245 1.225 8.245 0.45 3.435 0.45 3.435 1.225 3.205 1.225 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.285 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.17 0.515 3.17 0.515 3.75 0.285 3.75  ;
        POLYGON 4.065 1.28 4.61 1.28 4.61 1.51 4.295 1.51 4.295 3.685 4.065 3.685  ;
        POLYGON 2.325 1.315 2.715 1.315 2.715 3.055 3.735 3.055 3.735 3.975 5.755 3.975 5.755 4.315 3.505 4.315 3.505 3.285 2.555 3.285 2.555 3.685 2.325 3.685  ;
        POLYGON 6.105 3.045 8.375 3.045 8.375 3.855 8.145 3.855 8.145 3.275 6.335 3.275 6.335 3.855 6.105 3.855  ;
        POLYGON 5.085 2.765 5.445 2.765 5.445 1.225 5.675 1.225 5.675 2.585 9.59 2.585 9.59 2.815 5.67 2.815 5.67 2.995 5.315 2.995 5.315 3.685 5.085 3.685  ;
        POLYGON 6.67 1.95 9.635 1.95 9.635 1.225 9.865 1.225 9.865 2.13 10.115 2.13 10.115 3.995 9.885 3.995 9.885 2.36 9.64 2.36 9.64 2.18 6.67 2.18  ;
        POLYGON 6.125 1.455 9.175 1.455 9.175 0.765 11.575 0.765 11.575 3.065 11.345 3.065 11.345 0.995 10.55 0.995 10.55 2.025 10.32 2.025 10.32 0.995 9.405 0.995 9.405 1.685 6.355 1.685 6.355 2.025 6.125 2.025  ;
        POLYGON 11.9 1.225 12.155 1.225 12.155 3.525 11.9 3.525  ;
        POLYGON 10.78 1.225 11.01 1.225 11.01 3.185 11.135 3.185 11.135 3.765 14.72 3.765 14.72 2.725 14.95 2.725 14.95 3.995 10.78 3.995  ;
        POLYGON 12.58 2.725 12.81 2.725 12.81 3.295 14.26 3.295 14.26 2.265 15.44 2.265 15.44 1.315 15.67 1.315 15.67 1.975 15.93 1.975 15.93 2.495 14.49 2.495 14.49 3.525 12.58 3.525  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.6 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 1.77 3.895 1.77 3.895 2.15 2.945 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.38 1.675 14.41 1.675 14.41 2.15 13.38 2.15  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.575 1.77 1.575 2.245 0.71 2.245  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.51 3.45 17.685 3.45 17.685 0.845 17.915 0.845 17.915 3.83 17.51 3.83  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.225 4.59 3.225 3.045 3.455 3.045 3.455 4.59 5.99 4.59 7.305 4.59 7.305 3.515 7.535 3.515 7.535 4.59 8.555 4.59 9.045 4.59 9.045 3.44 9.275 3.44 9.275 4.59 9.77 4.59 10.295 4.59 13.525 4.59 13.525 4.345 13.755 4.345 13.755 4.59 15.495 4.59 15.845 4.59 15.845 3.875 16.075 3.875 16.075 4.59 16.665 4.59 16.665 3.875 16.895 3.875 16.895 4.59 17.39 4.59 18.705 4.59 18.705 3.875 18.935 3.875 18.935 4.59 19.6 4.59 19.6 5.49 17.39 5.49 15.495 5.49 10.295 5.49 9.77 5.49 8.555 5.49 5.99 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.6 -0.45 19.6 0.45 19.035 0.45 19.035 1.165 18.805 1.165 18.805 0.45 16.795 0.45 16.795 1.165 16.565 1.165 16.565 0.45 13.655 0.45 13.655 1.31 13.425 1.31 13.425 0.45 8.655 0.45 8.655 1.31 8.425 1.31 8.425 0.45 3.435 0.45 3.435 1.31 3.205 1.31 3.205 0.45 1.65 0.45 1.65 1.08 1.31 1.08 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.875 1.805 2.875 1.805 1.54 0.245 1.54 0.245 1.19 0.475 1.19 0.475 1.31 2.035 1.31 2.035 3.105 0.575 3.105 0.575 3.685 0.345 3.685  ;
        POLYGON 4.245 1.31 4.555 1.31 4.555 3.685 4.245 3.685  ;
        POLYGON 2.385 1.19 2.715 1.19 2.715 2.585 3.915 2.585 3.915 4.03 5.99 4.03 5.99 4.26 3.685 4.26 3.685 2.815 2.615 2.815 2.615 3.685 2.385 3.685  ;
        POLYGON 6.285 2.92 8.555 2.92 8.555 3.73 8.325 3.73 8.325 3.15 6.515 3.15 6.515 3.73 6.285 3.73  ;
        POLYGON 5.265 1.31 5.675 1.31 5.675 2.46 9.77 2.46 9.77 2.69 5.495 2.69 5.495 3.685 5.265 3.685  ;
        POLYGON 6.81 2 10.065 2 10.065 1.31 10.295 1.31 10.295 4.08 10.065 4.08 10.065 2.23 6.81 2.23  ;
        POLYGON 6.07 1.825 6.35 1.825 6.35 1.54 9.605 1.54 9.605 0.85 11.875 0.85 11.875 3.15 11.645 3.15 11.645 1.08 10.755 1.08 10.755 2.11 10.525 2.11 10.525 1.08 9.835 1.08 9.835 1.77 6.58 1.77 6.58 2.055 6.07 2.055  ;
        POLYGON 12.285 1.31 12.535 1.31 12.535 3.61 12.285 3.61  ;
        POLYGON 11.185 1.31 11.415 1.31 11.415 3.27 11.42 3.27 11.42 3.85 15.265 3.85 15.265 2.415 15.495 2.415 15.495 4.08 11.185 4.08  ;
        POLYGON 12.81 2.38 14.805 2.38 14.805 1.955 15.845 1.955 15.845 0.845 16.075 0.845 16.075 1.83 17.39 1.83 17.39 2.185 15.035 2.185 15.035 2.61 14.775 2.61 14.775 3.215 14.545 3.215 14.545 2.61 12.81 2.61  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.84 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.33 3.895 2.33 3.895 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.105 1.21 14.41 1.21 14.41 1.59 14.335 1.59 14.335 2.05 14.105 2.05  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.575 2.235 1.575 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.685 2.875 19.485 2.875 19.715 2.875 19.715 1.655 17.685 1.655 17.685 0.845 17.915 0.845 17.915 1.395 19.75 1.395 19.75 0.815 20.175 0.815 20.175 3.685 19.725 3.685 19.725 3.295 19.485 3.295 17.915 3.295 17.915 3.685 17.685 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.225 4.59 3.225 3.615 3.455 3.615 3.455 4.59 5.99 4.59 7.305 4.59 7.305 3.615 7.535 3.615 7.535 4.59 8.555 4.59 9.045 4.59 9.045 3.38 9.275 3.38 9.275 4.59 9.77 4.59 10.295 4.59 13.525 4.59 13.525 4.345 13.755 4.345 13.755 4.59 15.55 4.59 15.845 4.59 15.845 3.875 16.075 3.875 16.075 4.59 16.665 4.59 16.665 3.875 16.895 3.875 16.895 4.59 18.705 4.59 18.705 3.875 18.935 3.875 18.935 4.59 19.485 4.59 20.745 4.59 20.745 3.875 20.975 3.875 20.975 4.59 21.84 4.59 21.84 5.49 19.485 5.49 15.55 5.49 10.295 5.49 9.77 5.49 8.555 5.49 5.99 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.84 -0.45 21.84 0.45 21.275 0.45 21.275 1.165 21.045 1.165 21.045 0.45 19.035 0.45 19.035 1.165 18.805 1.165 18.805 0.45 16.795 0.45 16.795 1.165 16.565 1.165 16.565 0.45 13.655 0.45 13.655 1.25 13.425 1.25 13.425 0.45 8.955 0.45 8.955 1.25 8.725 1.25 8.725 0.45 3.435 0.45 3.435 1.25 3.205 1.25 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.245 1.25 4.555 1.25 4.555 3.785 4.245 3.785  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.155 3.915 3.155 3.915 4.13 5.99 4.13 5.99 4.36 3.685 4.36 3.685 3.385 2.615 3.385 2.615 3.685 2.385 3.685  ;
        POLYGON 6.285 3.145 8.555 3.145 8.555 3.955 8.325 3.955 8.325 3.375 6.515 3.375 6.515 3.955 6.285 3.955  ;
        POLYGON 5.265 1.25 5.675 1.25 5.675 2.685 9.77 2.685 9.77 2.915 5.495 2.915 5.495 3.785 5.265 3.785  ;
        POLYGON 6.81 2.225 10.065 2.225 10.065 1.25 10.295 1.25 10.295 4.02 10.065 4.02 10.065 2.455 6.81 2.455  ;
        POLYGON 6.07 1.765 9.605 1.765 9.605 0.79 11.875 0.79 11.875 3.09 11.645 3.09 11.645 1.02 10.755 1.02 10.755 2.05 10.525 2.05 10.525 1.02 9.835 1.02 9.835 1.995 6.07 1.995  ;
        POLYGON 12.285 1.25 12.535 1.25 12.535 3.55 12.285 3.55  ;
        POLYGON 11.185 1.25 11.415 1.25 11.415 3.21 11.42 3.21 11.42 3.79 15.07 3.79 15.07 2.47 15.55 2.47 15.55 2.7 15.3 2.7 15.3 4.02 11.185 4.02  ;
        POLYGON 12.81 2.32 14.61 2.32 14.61 2.01 15.845 2.01 15.845 0.845 16.075 0.845 16.075 2.015 19.485 2.015 19.485 2.275 15.845 2.275 15.845 2.24 14.84 2.24 14.84 3.215 14.555 3.215 14.555 2.55 12.81 2.55  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.33 3.975 2.33 3.975 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.965 2.2 17.77 2.2 17.77 2.76 16.965 2.76  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.545 2.33 15.575 2.33 15.575 2.805 14.545 2.805  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.575 2.235 1.575 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.685 0.845 20.01 0.845 20.01 3.685 19.705 3.685 19.705 1.655 19.685 1.655  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.515 3.535 3.515 3.535 4.59 7.605 4.59 7.605 4.375 7.835 4.375 7.835 4.59 10.805 4.59 10.805 4.375 11.035 4.375 11.035 4.59 12.715 4.59 14.85 4.59 14.85 3.95 15.19 3.95 15.19 4.59 16.89 4.59 16.89 3.95 17.23 3.95 17.23 4.59 18.69 4.59 18.985 4.59 18.985 3.425 19.215 3.425 19.215 4.59 19.475 4.59 20.725 4.59 20.725 3.875 20.955 3.875 20.955 4.59 21.28 4.59 21.28 5.49 19.475 5.49 18.69 5.49 12.715 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 21.035 0.45 21.035 1.165 20.805 1.165 20.805 0.45 17.175 0.45 17.175 1.225 16.945 1.225 16.945 0.45 9.175 0.45 9.175 1.425 8.945 1.425 8.945 0.45 3.435 0.45 3.435 1.425 3.205 1.425 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.655 1.315 0.655 1.51 2.035 1.51 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.325 1.315 4.555 1.315 4.555 3.685 4.325 3.685  ;
        POLYGON 6.365 3.345 9.075 3.345 9.075 3.685 6.365 3.685  ;
        POLYGON 5.345 2.685 5.825 2.685 5.825 1.315 6.055 1.315 6.055 2.685 10.005 2.685 10.005 2.575 10.235 2.575 10.235 2.915 5.575 2.915 5.575 3.685 5.345 3.685  ;
        POLYGON 9.565 3.345 11.39 3.345 11.39 2.345 7.335 2.345 7.335 2.455 7.105 2.455 7.105 2.115 11.425 2.115 11.425 1.315 11.655 1.315 11.655 3.445 12.045 3.445 12.045 2.875 12.275 2.875 12.275 3.685 9.565 3.685  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.055 3.995 3.055 3.995 3.915 12.715 3.915 12.715 4.315 12.485 4.315 12.485 4.145 6.07 4.145 6.07 4.26 3.765 4.26 3.765 3.285 2.615 3.285 2.615 3.685 2.385 3.685  ;
        POLYGON 6.285 1.655 10.965 1.655 10.965 0.68 14.555 0.68 14.555 1.64 14.325 1.64 14.325 0.91 11.195 0.91 11.195 1.885 6.515 1.885 6.515 2.115 6.285 2.115  ;
        POLYGON 13.665 1.315 13.895 1.315 13.895 1.87 14.985 1.87 14.985 1.315 15.215 1.315 15.215 1.87 16.155 1.87 16.155 3.215 15.925 3.215 15.925 2.1 14.315 2.1 14.315 3.215 14.085 3.215 14.085 2.115 13.665 2.115  ;
        POLYGON 12.545 1.315 13.295 1.315 13.295 3.455 18.46 3.455 18.46 2.415 18.69 2.415 18.69 3.685 13.065 3.685 13.065 1.655 12.545 1.655  ;
        POLYGON 17.965 2.885 18 2.885 18 1.97 16.735 1.97 16.735 2.115 16.505 2.115 16.505 1.74 18.905 1.74 18.905 1.315 19.135 1.315 19.135 1.975 19.475 1.975 19.475 2.315 18.91 2.315 18.91 2.025 18.23 2.025 18.23 3.225 17.965 3.225  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 22.4 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.39 1.77 3.99 1.77 3.99 1.21 4.33 1.21 4.33 2.15 3.39 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.755 2.32 17.77 2.32 17.77 2.71 16.755 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.27 1.21 15.61 1.21 15.61 2.06 15.27 2.06  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.58 1.77 1.58 2.15 0.71 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.67 0.845 21.13 0.845 21.13 3.83 20.67 3.83  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.47 4.59 1.47 3.425 1.7 3.425 1.7 4.59 2.14 4.59 3.21 4.59 3.21 3.595 3.44 3.595 3.44 4.59 7.69 4.59 7.69 4.48 7.92 4.48 7.92 4.59 10.83 4.59 10.83 4.48 11.06 4.48 11.06 4.59 12.795 4.59 14.775 4.59 14.775 3.96 15.115 3.96 15.115 4.59 16.815 4.59 16.815 3.96 17.155 3.96 17.155 4.59 18.69 4.59 18.91 4.59 18.91 3.905 19.14 3.905 19.14 4.59 19.65 4.59 19.65 3.875 19.88 3.875 19.88 4.59 20.32 4.59 21.69 4.59 21.69 3.875 21.92 3.875 21.92 4.59 22.4 4.59 22.4 5.49 20.32 5.49 18.69 5.49 12.795 5.49 2.14 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 22.4 -0.45 22.4 0.45 22.02 0.45 22.02 1.165 21.79 1.165 21.79 0.45 19.78 0.45 19.78 1.165 19.55 1.165 19.55 0.45 17.1 0.45 17.1 1.225 16.87 1.225 16.87 0.45 9.215 0.45 9.215 1.37 8.875 1.37 8.875 0.45 3.67 0.45 3.67 1.425 3.44 1.425 3.44 0.45 1.755 0.45 1.755 1.045 1.415 1.045 1.415 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.45 2.875 1.91 2.875 1.91 1.54 0.35 1.54 0.35 1.19 0.58 1.19 0.58 1.31 2.14 1.31 2.14 3.105 0.68 3.105 0.68 3.685 0.45 3.685  ;
        POLYGON 4.23 2.955 4.56 2.955 4.56 1.315 4.79 1.315 4.79 3.185 4.46 3.185 4.46 3.765 4.23 3.765  ;
        POLYGON 6.52 2.98 6.75 2.98 6.75 3.45 9.16 3.45 9.16 3.79 6.52 3.79  ;
        POLYGON 5.25 2.52 5.68 2.52 5.68 1.315 5.91 1.315 5.91 2.52 10.09 2.52 10.09 2.505 10.32 2.505 10.32 2.845 10.09 2.845 10.09 2.75 5.48 2.75 5.48 3.765 5.25 3.765  ;
        POLYGON 9.65 2.98 9.88 2.98 9.88 3.075 10.55 3.075 10.55 2.275 10.005 2.275 10.005 2.29 7.1 2.29 7.1 1.95 7.33 1.95 7.33 2.06 9.92 2.06 9.92 2.045 11.21 2.045 11.21 1.315 11.44 1.315 11.44 2.225 12.3 2.225 12.3 3.775 12.07 3.775 12.07 2.455 10.78 2.455 10.78 3.305 9.88 3.305 9.88 3.79 9.65 3.79  ;
        POLYGON 2.49 1.19 2.82 1.19 2.82 2.985 3.9 2.985 3.9 4.02 12.795 4.02 12.795 4.35 12.455 4.35 12.455 4.25 5.975 4.25 5.975 4.34 3.67 4.34 3.67 3.215 2.49 3.215  ;
        POLYGON 6.36 1.49 7.73 1.49 7.73 1.6 9.605 1.6 9.605 0.68 14.38 0.68 14.38 0.91 9.835 0.91 9.835 1.83 7.53 1.83 7.53 1.72 6.59 1.72 6.59 2.115 6.36 2.115  ;
        POLYGON 13.45 1.14 14.81 1.14 14.81 0.75 16.08 0.75 16.08 3.225 15.85 3.225 15.85 0.98 15.04 0.98 15.04 1.37 14.34 1.37 14.34 3.305 14.11 3.305 14.11 1.48 13.45 1.48  ;
        POLYGON 12.33 1.315 12.56 1.315 12.56 1.67 13.32 1.67 13.32 3.545 14.495 3.545 14.495 3.5 18.46 3.5 18.46 2.425 18.69 2.425 18.69 3.73 14.635 3.73 14.635 3.775 13.09 3.775 13.09 1.9 12.33 1.9  ;
        POLYGON 17.89 2.91 18 2.91 18 2.09 16.375 2.09 16.375 1.86 18.83 1.86 18.83 1.315 19.06 1.315 19.06 1.775 20.32 1.775 20.32 2.115 18.23 2.115 18.23 3.25 17.89 3.25  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.64 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.055 2.33 3.89 2.33 3.89 2.71 3.055 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.95 2.48 17.515 2.48 17.515 2.71 17.21 2.71 17.21 3.27 16.95 3.27  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.27 1.77 15.53 1.77 15.53 2.765 15.27 2.765  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.295 1.57 2.295 1.57 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.59 2.875 22.435 2.875 22.665 2.875 22.665 1.655 20.59 1.655 20.59 0.845 20.82 0.845 20.82 1.395 22.55 1.395 22.55 0.815 23.06 0.815 23.06 3.685 22.63 3.685 22.63 3.105 22.435 3.105 20.82 3.105 20.82 3.685 20.59 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.205 4.59 3.205 3.515 3.435 3.515 3.435 4.59 7.465 4.59 7.465 4.49 7.695 4.49 7.695 4.59 10.665 4.59 10.665 4.49 10.895 4.49 10.895 4.59 12.63 4.59 14.695 4.59 14.695 3.96 15.035 3.96 15.035 4.59 16.735 4.59 16.735 3.96 17.075 3.96 17.075 4.59 18.5 4.59 18.83 4.59 18.83 3.435 19.06 3.435 19.06 4.59 19.57 4.59 19.57 3.875 19.8 3.875 19.8 4.59 21.61 4.59 21.61 3.875 21.84 3.875 21.84 4.59 22.435 4.59 23.65 4.59 23.65 3.875 23.88 3.875 23.88 4.59 24.64 4.59 24.64 5.49 22.435 5.49 18.5 5.49 12.63 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 24.64 -0.45 24.64 0.45 24.18 0.45 24.18 1.165 23.95 1.165 23.95 0.45 21.94 0.45 21.94 1.165 21.71 1.165 21.71 0.45 19.7 0.45 19.7 1.165 19.47 1.165 19.47 0.45 17.02 0.45 17.02 1.225 16.79 1.225 16.79 0.45 8.635 0.45 8.635 1.425 8.405 1.425 8.405 0.45 3.435 0.45 3.435 1.425 3.205 1.425 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.225 1.315 4.555 1.315 4.555 3.685 4.225 3.685  ;
        POLYGON 6.285 3.35 8.935 3.35 8.935 3.8 6.285 3.8  ;
        POLYGON 5.245 1.315 5.675 1.315 5.675 2.685 9.865 2.685 9.865 2.575 10.095 2.575 10.095 2.915 5.475 2.915 5.475 3.685 5.245 3.685  ;
        POLYGON 9.425 3.46 11.285 3.46 11.285 2.345 7.095 2.345 7.095 2.455 6.865 2.455 6.865 2.115 11.285 2.115 11.285 1.315 11.515 1.315 11.515 3.57 11.905 3.57 11.905 2.875 12.135 2.875 12.135 3.8 9.425 3.8  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.055 3.895 3.055 3.895 4.03 12.63 4.03 12.63 4.26 3.665 4.26 3.665 3.285 2.615 3.285 2.615 3.685 2.385 3.685  ;
        POLYGON 6.125 1.655 10.825 1.655 10.825 0.68 14.455 0.68 14.455 0.91 11.055 0.91 11.055 1.885 6.355 1.885 6.355 2.115 6.125 2.115  ;
        POLYGON 13.525 1.31 16 1.31 16 3.225 15.77 3.225 15.77 1.54 14.175 1.54 14.175 3.215 13.945 3.215 13.945 1.655 13.525 1.655  ;
        POLYGON 12.405 1.315 13.155 1.315 13.155 3.5 18.27 3.5 18.27 2.425 18.5 2.425 18.5 3.73 12.925 3.73 12.925 1.655 12.405 1.655  ;
        POLYGON 16.295 1.83 18.75 1.83 18.75 1.315 18.98 1.315 18.98 1.775 20.24 1.775 20.24 2.005 22.435 2.005 22.435 2.29 20.01 2.29 20.01 2.115 18.04 2.115 18.04 3.225 17.81 3.225 17.81 2.06 16.295 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.16 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 2.33 4.55 2.33 4.55 2.71 3.51 2.71  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.15 2.265 14.975 2.265 14.975 2.71 14.15 2.71  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.77 1.53 1.77 1.53 2.15 0.63 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.07 0.845 18.375 0.845 18.375 3.685 18.145 3.685 18.145 1.59 18.07 1.59  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.425 1.495 3.425 1.495 4.59 2.035 4.59 3.005 4.59 3.005 3.905 3.235 3.905 3.235 4.59 7.245 4.59 7.245 3.905 7.475 3.905 7.475 4.59 9.725 4.59 9.725 3.905 9.955 3.905 9.955 4.59 11.535 4.59 13.805 4.59 13.805 3.915 14.035 3.915 14.035 4.59 16.345 4.59 16.345 3.175 16.575 3.175 16.575 4.59 17.07 4.59 17.915 4.59 19.165 4.59 19.165 3.875 19.395 3.875 19.395 4.59 20.16 4.59 20.16 5.49 17.915 5.49 17.07 5.49 11.535 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.16 -0.45 20.16 0.45 19.495 0.45 19.495 1.165 19.265 1.165 19.265 0.45 16.535 0.45 16.535 1.42 16.305 1.42 16.305 0.45 7.655 0.45 7.655 1.425 7.425 1.425 7.425 0.45 3.455 0.45 3.455 1.425 3.225 1.425 3.225 0.45 1.595 0.45 1.595 1.08 1.365 1.08 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.875 1.805 2.875 1.805 1.54 0.245 1.54 0.245 1.17 0.475 1.17 0.475 1.31 2.035 1.31 2.035 3.105 0.475 3.105 0.475 3.685 0.245 3.685  ;
        POLYGON 3.05 1.87 3.685 1.87 3.685 1.315 4.575 1.315 4.575 1.655 3.915 1.655 3.915 2.1 3.28 2.1 3.28 2.985 4.53 2.985 4.53 3.215 3.05 3.215  ;
        POLYGON 5.265 1.315 5.695 1.315 5.695 1.83 8.19 1.83 8.19 2.06 5.495 2.06 5.495 3.215 5.265 3.215  ;
        POLYGON 6.53 2.47 9.425 2.47 9.425 1.315 9.655 1.315 9.655 2.47 11.095 2.47 11.095 3.215 10.865 3.215 10.865 2.7 8.715 2.7 8.715 3.215 8.485 3.215 8.485 2.7 6.53 2.7  ;
        POLYGON 2.285 1.17 2.715 1.17 2.715 3.445 11.535 3.445 11.535 4.315 11.305 4.315 11.305 3.675 5.99 3.675 5.99 4.26 5.65 4.26 5.65 3.675 2.515 3.675 2.515 3.685 2.285 3.685  ;
        POLYGON 13.085 2.875 13.69 2.875 13.69 1.545 11.845 1.545 11.845 1.205 13.92 1.205 13.92 2.985 15.105 2.985 15.105 2.905 15.335 2.905 15.335 3.245 15.105 3.245 15.105 3.215 13.085 3.215  ;
        POLYGON 10.725 1.315 10.955 1.315 10.955 1.775 12.115 1.775 12.115 3.455 14.225 3.455 14.225 3.475 15.885 3.475 15.885 2.5 17.07 2.5 17.07 2.73 16.115 2.73 16.115 3.705 14.13 3.705 14.13 3.685 11.885 3.685 11.885 2.005 10.725 2.005  ;
        POLYGON 15.685 1.93 17.425 1.93 17.425 1.315 17.655 1.315 17.655 1.975 17.915 1.975 17.915 2.315 17.595 2.315 17.595 3.715 17.365 3.715 17.365 2.27 15.685 2.27  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.83 1.96 4.63 1.96 4.63 1.77 4.89 1.77 4.89 2.19 3.83 2.19  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.655 2.165 14.86 2.165 14.86 2.71 13.655 2.71  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.575 2.235 1.575 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.12 0.845 19.45 0.845 19.45 3.685 19.12 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.58 3.535 3.58 3.535 4.59 7.305 4.59 7.305 3.11 7.535 3.11 7.535 4.59 9.365 4.59 9.365 3.11 9.595 3.11 9.595 4.59 11.435 4.59 13.745 4.59 13.745 3.97 13.975 3.97 13.975 4.59 16.345 4.59 16.345 3.21 16.575 3.21 16.575 4.59 17.07 4.59 18.1 4.59 18.1 3.875 18.33 3.875 18.33 4.59 18.77 4.59 20.14 4.59 20.14 3.875 20.37 3.875 20.37 4.59 21.28 4.59 21.28 5.49 18.77 5.49 17.07 5.49 11.435 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.57 0.45 20.57 1.165 20.34 1.165 20.34 0.45 18.33 0.45 18.33 1.165 18.1 1.165 18.1 0.45 16.475 0.45 16.475 1.42 16.245 1.42 16.245 0.45 7.635 0.45 7.635 1.325 7.405 1.325 7.405 0.45 3.49 0.45 3.49 1.27 3.15 1.27 3.15 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.9 0.575 2.9 0.575 2.94 1.805 2.94 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.17 0.575 3.17 0.575 3.71 0.345 3.71  ;
        POLYGON 3.6 2.42 4.555 2.42 4.555 3.75 4.325 3.75 4.325 2.65 3.37 2.65 3.37 1.5 3.715 1.5 3.715 1.32 4.325 1.32 4.325 1.21 4.555 1.21 4.555 1.55 3.94 1.55 3.94 1.73 3.6 1.73  ;
        POLYGON 5.445 1.215 5.675 1.215 5.675 1.73 8.13 1.73 8.13 1.96 5.675 1.96 5.675 3.75 5.445 3.75  ;
        POLYGON 6.81 2.19 9.365 2.19 9.365 1.215 9.595 1.215 9.595 2.19 10.995 2.19 10.995 3.685 10.765 3.685 10.765 2.42 8.555 2.42 8.555 3.75 8.325 3.75 8.325 2.42 6.81 2.42  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 2.985 3.995 2.985 3.995 4.095 6.845 4.095 6.845 2.65 7.995 2.65 7.995 3.98 8.905 3.98 8.905 2.65 10.055 2.65 10.055 3.975 11.435 3.975 11.435 4.315 9.825 4.315 9.825 2.88 9.135 2.88 9.135 4.21 7.765 4.21 7.765 2.88 7.075 2.88 7.075 4.325 3.765 4.325 3.765 3.215 2.385 3.215  ;
        POLYGON 13.255 2.94 15.275 2.94 15.275 3.28 13.025 3.28 13.025 1.5 11.785 1.5 11.785 1.16 13.875 1.16 13.875 1.5 13.255 1.5  ;
        POLYGON 10.665 1.215 10.895 1.215 10.895 1.73 12.015 1.73 12.015 3.51 15.885 3.51 15.885 2.535 17.07 2.535 17.07 2.765 16.115 2.765 16.115 3.74 11.785 3.74 11.785 1.96 10.665 1.96  ;
        POLYGON 15.625 1.775 17.365 1.775 17.365 1.315 17.595 1.315 17.595 1.775 18.77 1.775 18.77 2.115 17.595 2.115 17.595 3.75 17.365 3.75 17.365 2.115 15.625 2.115  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 2.33 4.525 2.33 4.525 2.71 3.51 2.71  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 2.15 15.53 2.15 15.53 2.71 14.71 2.71  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.24 1.575 2.24 1.575 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.665 2.875 21.425 2.875 21.655 2.875 21.655 1.655 19.665 1.655 19.665 0.845 19.895 0.845 19.895 1.395 21.43 1.395 21.43 0.815 22.135 0.815 22.135 3.685 21.705 3.685 21.705 3.105 21.425 3.105 19.895 3.105 19.895 3.685 19.665 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.105 4.59 3.105 3.86 3.335 3.86 3.335 4.59 7.345 4.59 7.345 3.905 7.575 3.905 7.575 4.59 9.825 4.59 9.825 3.905 10.055 3.905 10.055 4.59 11.795 4.59 14.205 4.59 14.205 3.915 14.435 3.915 14.435 4.59 16.745 4.59 16.745 3.155 16.975 3.155 16.975 4.59 17.47 4.59 18.645 4.59 18.645 3.875 18.875 3.875 18.875 4.59 20.685 4.59 20.685 3.875 20.915 3.875 20.915 4.59 21.425 4.59 22.725 4.59 22.725 3.875 22.955 3.875 22.955 4.59 23.52 4.59 23.52 5.49 21.425 5.49 17.47 5.49 11.795 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 23.255 0.45 23.255 1.165 23.025 1.165 23.025 0.45 21.015 0.45 21.015 1.165 20.785 1.165 20.785 0.45 18.775 0.45 18.775 1.165 18.545 1.165 18.545 0.45 16.755 0.45 16.755 1.425 16.525 1.425 16.525 0.45 7.755 0.45 7.755 1.425 7.525 1.425 7.525 0.45 3.455 0.45 3.455 1.425 3.225 1.425 3.225 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 1.685 0.245 1.685 0.245 1.315 0.475 1.315 0.475 1.455 2.035 1.455 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 3.28 2.94 4.63 2.94 4.63 3.205 4.29 3.205 4.29 3.17 3.05 3.17 3.05 1.87 4.345 1.87 4.345 1.315 4.575 1.315 4.575 2.1 3.28 2.1  ;
        POLYGON 5.365 1.315 5.795 1.315 5.795 1.83 8.29 1.83 8.29 2.06 5.595 2.06 5.595 3.26 5.365 3.26  ;
        POLYGON 6.63 2.515 9.825 2.515 9.825 1.315 10.055 1.315 10.055 2.515 11.355 2.515 11.355 3.215 11.125 3.215 11.125 2.745 8.815 2.745 8.815 3.215 8.585 3.215 8.585 2.745 6.63 2.745  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.4 3.705 3.4 3.705 3.49 5.895 3.49 5.895 3.445 11.795 3.445 11.795 4.315 11.565 4.315 11.565 3.675 6.035 3.675 6.035 4.36 5.805 4.36 5.805 3.72 3.52 3.72 3.52 3.63 2.615 3.63 2.615 3.685 2.385 3.685  ;
        POLYGON 13.485 2.875 14.105 2.875 14.105 1.545 12.245 1.545 12.245 1.205 14.335 1.205 14.335 2.995 15.79 2.995 15.79 3.225 13.485 3.225  ;
        POLYGON 11.125 1.315 11.355 1.315 11.355 1.775 12.375 1.775 12.375 3.455 16.285 3.455 16.285 2.48 17.47 2.48 17.47 2.71 16.515 2.71 16.515 3.685 12.145 3.685 12.145 2.005 11.125 2.005  ;
        POLYGON 16.085 1.775 17.825 1.775 17.825 1.315 18.055 1.315 18.055 1.96 21.425 1.96 21.425 2.32 17.995 2.32 17.995 3.695 17.765 3.695 17.765 2.115 16.085 2.115  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.21 4.89 1.21 4.89 2.115 4.63 2.115  ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.575 2.235 1.575 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 2.33 14.885 2.33 14.885 0.845 15.115 0.845 15.115 3.685 14.71 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.895 1.595 3.895 1.595 4.59 3.185 4.59 3.185 3.905 3.415 3.905 3.415 4.59 6.115 4.59 7.205 4.59 7.205 3.045 7.435 3.045 7.435 4.59 7.875 4.59 8.855 4.59 12.025 4.59 12.025 3.145 12.255 3.145 12.255 4.59 12.75 4.59 13.765 4.59 13.765 3.875 13.995 3.875 13.995 4.59 14.49 4.59 15.68 4.59 15.68 5.49 14.49 5.49 12.75 5.49 8.855 5.49 7.875 5.49 6.115 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 13.995 0.45 13.995 1.165 13.765 1.165 13.765 0.45 12.155 0.45 12.155 1.265 11.925 1.265 11.925 0.45 7.525 0.45 7.525 0.625 7.295 0.625 7.295 0.45 3.435 0.45 3.435 1.435 3.205 1.435 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 3.425 1.805 3.425 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.445 6.115 3.445 6.115 4.315 5.885 4.315 5.885 3.675 1.94 3.675 1.94 3.655 0.575 3.655 0.575 4.235 0.345 4.235  ;
        POLYGON 5.165 1.315 5.395 1.315 5.395 2.415 7.875 2.415 7.875 2.755 5.395 2.755 5.395 3.215 5.165 3.215  ;
        POLYGON 6.685 1.775 8.225 1.775 8.225 1.315 8.855 1.315 8.855 1.655 8.455 1.655 8.455 3.685 8.225 3.685 8.225 2.115 6.685 2.115  ;
        POLYGON 2.385 2.525 3.845 2.525 3.845 1.895 2.485 1.895 2.485 1.315 2.715 1.315 2.715 1.665 3.845 1.665 3.845 0.69 5.89 0.69 5.89 0.855 9.01 0.855 9.01 0.69 10.735 0.69 10.735 2.755 10.505 2.755 10.505 1.085 5.665 1.085 5.665 0.92 4.075 0.92 4.075 2.755 2.615 2.755 2.615 3.215 2.385 3.215  ;
        POLYGON 9.745 1.315 9.975 1.315 9.975 3.455 11.565 3.455 11.565 2.47 12.75 2.47 12.75 2.7 11.795 2.7 11.795 3.685 9.745 3.685  ;
        POLYGON 11.265 1.775 13.045 1.775 13.045 1.315 13.275 1.315 13.275 1.83 14.49 1.83 14.49 2.06 13.275 2.06 13.275 3.685 13.045 3.685 13.045 2.115 11.265 2.115  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 16.8 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.21 5.08 1.21 5.08 2.05 4.63 2.05  ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.77 1.49 1.77 1.49 2.15 0.63 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 1.21 15.095 1.21 15.095 0.845 15.325 0.845 15.325 3.685 14.995 3.685 14.995 1.59 14.71 1.59  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.21 4.59 1.21 3.95 1.55 3.95 1.55 4.59 3.395 4.59 3.395 3.885 3.625 3.885 3.625 4.59 6.145 4.59 7.235 4.59 7.235 3.09 7.465 3.09 7.465 4.59 8.085 4.59 9.065 4.59 12.235 4.59 12.235 3.875 12.465 3.875 12.465 4.59 12.96 4.59 13.975 4.59 13.975 3.875 14.205 3.875 14.205 4.59 14.7 4.59 16.015 4.59 16.015 3.875 16.245 3.875 16.245 4.59 16.8 4.59 16.8 5.49 14.7 5.49 12.96 5.49 9.065 5.49 8.085 5.49 6.145 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 16.8 -0.45 16.8 0.45 16.445 0.45 16.445 1.165 16.215 1.165 16.215 0.45 14.205 0.45 14.205 1.165 13.975 1.165 13.975 0.45 12.365 0.45 12.365 1.16 12.135 1.16 12.135 0.45 7.785 0.45 7.785 0.545 7.555 0.545 7.555 0.45 3.425 0.45 3.425 0.665 1.595 0.665 1.595 1.08 1.365 1.08 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.425 1.805 3.425 1.805 1.54 0.245 1.54 0.245 1.17 0.475 1.17 0.475 1.31 2.035 1.31 2.035 3.445 3.205 3.445 3.205 3.425 4.085 3.425 4.085 4.02 6.145 4.02 6.145 4.36 3.855 4.36 3.855 3.655 3.3 3.655 3.3 3.675 0.475 3.675 0.475 4.235 0.245 4.235  ;
        POLYGON 5.375 1.305 5.605 1.305 5.605 2.46 8.085 2.46 8.085 2.8 5.605 2.8 5.605 3.73 5.375 3.73  ;
        POLYGON 6.655 1.765 8.835 1.765 8.835 1.31 9.065 1.31 9.065 3.73 8.835 3.73 8.835 2.105 6.655 2.105  ;
        POLYGON 2.385 1.17 2.715 1.17 2.715 2.57 4.055 2.57 4.055 0.68 6.1 0.68 6.1 0.775 9.22 0.775 9.22 0.685 10.945 0.685 10.945 2.8 10.715 2.8 10.715 1.005 5.995 1.005 5.995 0.98 4.285 0.98 4.285 2.8 2.615 2.8 2.615 3.215 2.385 3.215  ;
        POLYGON 9.955 1.31 10.185 1.31 10.185 3.5 11.825 3.5 11.825 2.47 12.96 2.47 12.96 2.7 12.055 2.7 12.055 3.73 9.955 3.73  ;
        POLYGON 11.475 1.77 13.255 1.77 13.255 0.84 13.485 0.84 13.485 1.83 14.7 1.83 14.7 2.06 13.485 2.06 13.485 3.685 13.255 3.685 13.255 2.11 11.475 2.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.6 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.21 4.89 1.21 4.89 2.115 4.63 2.115  ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.505 2.235 1.505 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.125 2.875 16.885 2.875 17.115 2.875 17.115 1.655 15.285 1.655 15.285 0.845 15.515 0.845 15.515 1.395 17.51 1.395 17.51 0.815 17.77 0.815 17.77 3.685 17.165 3.685 17.165 3.105 16.885 3.105 15.355 3.105 15.355 3.685 15.125 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.31 4.59 1.31 3.95 1.65 3.95 1.65 4.59 3.185 4.59 3.185 3.905 3.415 3.905 3.415 4.59 6.035 4.59 7.125 4.59 7.125 3.045 7.355 3.045 7.355 4.59 8.175 4.59 8.855 4.59 12.065 4.59 12.065 3.875 12.295 3.875 12.295 4.59 12.79 4.59 14.105 4.59 14.105 3.875 14.335 3.875 14.335 4.59 16.145 4.59 16.145 3.875 16.375 3.875 16.375 4.59 16.885 4.59 18.185 4.59 18.185 3.875 18.415 3.875 18.415 4.59 19.6 4.59 19.6 5.49 16.885 5.49 12.79 5.49 8.855 5.49 8.175 5.49 6.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.6 -0.45 19.6 0.45 18.875 0.45 18.875 1.165 18.645 1.165 18.645 0.45 16.635 0.45 16.635 1.165 16.405 1.165 16.405 0.45 14.395 0.45 14.395 1.165 14.165 1.165 14.165 0.45 12.155 0.45 12.155 1.165 11.925 1.165 11.925 0.45 7.52 0.45 7.52 0.625 7.29 0.625 7.29 0.45 3.435 0.45 3.435 1.435 3.205 1.435 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 3.425 1.805 3.425 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.445 6.035 3.445 6.035 4.315 5.805 4.315 5.805 3.675 0.575 3.675 0.575 4.235 0.345 4.235  ;
        POLYGON 5.165 1.315 5.395 1.315 5.395 2.415 8.175 2.415 8.175 2.755 5.395 2.755 5.395 3.215 5.165 3.215  ;
        POLYGON 6.685 1.775 8.625 1.775 8.625 1.315 8.855 1.315 8.855 3.685 8.62 3.685 8.62 2.115 6.685 2.115  ;
        POLYGON 2.385 2.525 3.845 2.525 3.845 1.895 2.485 1.895 2.485 1.315 2.715 1.315 2.715 1.665 3.845 1.665 3.845 0.69 5.89 0.69 5.89 0.855 9.01 0.855 9.01 0.69 10.855 0.69 10.855 2.755 10.625 2.755 10.625 1.085 5.665 1.085 5.665 0.92 4.075 0.92 4.075 2.755 2.615 2.755 2.615 3.215 2.385 3.215  ;
        POLYGON 9.745 1.315 9.975 1.315 9.975 3.455 11.705 3.455 11.705 2.47 12.79 2.47 12.79 2.7 11.935 2.7 11.935 3.685 9.745 3.685  ;
        POLYGON 11.265 1.775 13.045 1.775 13.045 0.845 13.31 0.845 13.31 1.975 16.885 1.975 16.885 2.315 13.315 2.315 13.315 3.685 13.085 3.685 13.085 2.115 11.265 2.115  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.28 2.33 3.915 2.33 3.915 2.71 3.28 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.83 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.865 1.66 14.15 1.66 14.15 1.21 15.07 1.21 15.07 1.59 14.38 1.59 14.38 2 13.865 2  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 2.15 0.97 2.15 0.97 2.71 0.66 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.325 0.845 16.65 0.845 16.65 3.685 16.345 3.685 16.345 2.19 16.325 2.19  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.285 4.59 1.285 3.425 1.515 3.425 1.515 4.59 2.01 4.59 3.245 4.59 3.245 3.615 3.475 3.615 3.475 4.59 4.99 4.59 7.325 4.59 7.325 3.615 7.555 3.615 7.555 4.59 8.575 4.59 9.065 4.59 9.065 3.33 9.295 3.33 9.295 4.59 9.79 4.59 10.315 4.59 13.365 4.59 13.365 4.19 13.595 4.19 13.595 4.59 15.295 4.59 15.625 4.59 15.625 3.31 15.855 3.31 15.855 4.59 16.1 4.59 17.365 4.59 17.365 3.875 17.595 3.875 17.595 4.59 17.92 4.59 17.92 5.49 16.1 5.49 15.295 5.49 10.315 5.49 9.79 5.49 8.575 5.49 4.99 5.49 2.01 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.675 0.45 17.675 1.165 17.445 1.165 17.445 0.45 13.415 0.45 13.415 1.2 13.185 1.2 13.185 0.45 8.935 0.45 8.935 1.2 8.705 1.2 8.705 0.45 3.455 0.45 3.455 1.2 3.225 1.2 3.225 0.45 1.615 0.45 1.615 1.225 1.385 1.225 1.385 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.265 2.875 0.495 2.875 0.495 2.94 1.2 2.94 1.2 1.685 0.21 1.685 0.21 1.37 1.085 1.37 1.085 1.455 1.43 1.455 1.43 2.03 2.01 2.03 2.01 2.26 1.43 2.26 1.43 3.17 0.495 3.17 0.495 3.685 0.265 3.685  ;
        POLYGON 4.265 1.2 4.575 1.2 4.575 3.785 4.265 3.785  ;
        POLYGON 2.305 1.315 2.735 1.315 2.735 3.155 3.935 3.155 3.935 4.13 4.99 4.13 4.99 4.36 3.705 4.36 3.705 3.385 2.535 3.385 2.535 3.685 2.305 3.685  ;
        POLYGON 6.305 3.145 8.575 3.145 8.575 3.955 8.345 3.955 8.345 3.375 6.535 3.375 6.535 3.955 6.305 3.955  ;
        POLYGON 5.52 2.685 9.79 2.685 9.79 2.915 5.515 2.915 5.515 3.785 5.285 3.785 5.285 1.2 5.695 1.2 5.695 1.54 5.52 1.54  ;
        POLYGON 6.83 2.175 9.825 2.175 9.825 1.2 10.055 1.2 10.055 2.23 10.315 2.23 10.315 3.97 10.085 3.97 10.085 2.46 9.855 2.46 9.855 2.405 6.83 2.405  ;
        POLYGON 5.85 1.715 9.365 1.715 9.365 0.74 11.83 0.74 11.83 2.985 11.485 2.985 11.485 0.97 10.515 0.97 10.515 2 10.285 2 10.285 0.97 9.595 0.97 9.595 1.945 5.85 1.945  ;
        POLYGON 12.065 1.2 12.355 1.2 12.355 3.5 12.065 3.5  ;
        POLYGON 10.945 1.2 11.175 1.2 11.175 3.16 11.335 3.16 11.335 3.73 15.065 3.73 15.065 2.7 15.295 2.7 15.295 3.96 11.335 3.96 11.335 3.97 10.945 3.97  ;
        POLYGON 12.65 2.24 15.605 2.24 15.605 1.29 15.835 1.29 15.835 2.24 16.1 2.24 16.1 2.47 14.835 2.47 14.835 3.5 14.605 3.5 14.605 2.65 12.65 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.96 2.33 3.895 2.33 3.895 2.71 2.96 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.59 2.33 14.015 2.33 14.015 2.71 13.59 2.71  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.265 1.59 2.265 1.59 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6016 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.445 0.845 17.77 0.845 17.77 3.685 17.445 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.09 4.59 3.225 4.59 3.225 3.615 3.455 3.615 3.455 4.59 4.97 4.59 7.305 4.59 7.305 3.615 7.535 3.615 7.535 4.59 8.555 4.59 9.045 4.59 9.045 3.32 9.275 3.32 9.275 4.59 9.77 4.59 10.295 4.59 13.345 4.59 13.345 4.345 13.575 4.345 13.575 4.59 15.155 4.59 15.385 4.59 15.385 3.875 15.615 3.875 15.615 4.59 16.425 4.59 16.425 3.875 16.655 3.875 16.655 4.59 17.05 4.59 18.465 4.59 18.465 3.875 18.695 3.875 18.695 4.59 19.04 4.59 19.04 5.49 17.05 5.49 15.155 5.49 10.295 5.49 9.77 5.49 8.555 5.49 4.97 5.49 2.09 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 18.795 0.45 18.795 1.235 18.565 1.235 18.565 0.45 16.555 0.45 16.555 1.235 16.325 1.235 16.325 0.45 13.365 0.45 13.365 1.195 13.135 1.195 13.135 0.45 8.655 0.45 8.655 1.195 8.425 1.195 8.425 0.45 3.435 0.45 3.435 1.195 3.205 1.195 3.205 0.45 1.595 0.45 1.595 1.2 1.365 1.2 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.925 0.575 2.925 0.575 2.965 1.86 2.965 1.86 2.035 0.245 2.035 0.245 1.29 0.475 1.29 0.475 1.805 2.09 1.805 2.09 3.195 0.575 3.195 0.575 3.735 0.345 3.735  ;
        POLYGON 4.245 1.195 4.555 1.195 4.555 3.785 4.245 3.785  ;
        POLYGON 2.385 1.29 2.715 1.29 2.715 3.155 3.915 3.155 3.915 4.13 4.97 4.13 4.97 4.36 3.685 4.36 3.685 3.385 2.615 3.385 2.615 3.685 2.385 3.685  ;
        POLYGON 6.285 3.145 8.555 3.145 8.555 3.955 8.325 3.955 8.325 3.375 6.515 3.375 6.515 3.955 6.285 3.955  ;
        POLYGON 5.495 2.685 9.77 2.685 9.77 2.915 5.495 2.915 5.495 3.785 5.265 3.785 5.265 1.185 5.675 1.185 5.675 1.525 5.495 1.525  ;
        POLYGON 6.81 2.225 9.765 2.225 9.765 1.195 9.995 1.195 9.995 2.225 10.295 2.225 10.295 3.96 10.065 3.96 10.065 2.455 6.81 2.455  ;
        POLYGON 5.855 1.71 9.305 1.71 9.305 0.735 11.785 0.735 11.785 2.69 11.815 2.69 11.815 3.03 11.555 3.03 11.555 0.965 10.455 0.965 10.455 1.995 10.225 1.995 10.225 0.965 9.535 0.965 9.535 1.94 5.855 1.94  ;
        POLYGON 12.015 1.195 12.335 1.195 12.335 3.49 12.105 3.49 12.105 1.535 12.015 1.535  ;
        POLYGON 10.895 1.195 11.315 1.195 11.315 3.73 14.925 3.73 14.925 2.415 15.155 2.415 15.155 3.96 10.895 3.96  ;
        POLYGON 12.63 2.745 12.97 2.745 12.97 2.94 14.465 2.94 14.465 1.955 15.555 1.955 15.555 0.725 15.785 0.725 15.785 1.83 17.05 1.83 17.05 2.185 14.695 2.185 14.695 3.17 12.63 3.17  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.75 3.895 1.75 3.895 2.09 2.89 2.09  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.97 1.75 13.78 1.75 13.78 2.09 12.97 2.09  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.33 1.57 2.33 1.57 2.71 0.15 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.37 2.875 19.365 2.875 19.595 2.875 19.595 1.625 17.37 1.625 17.37 0.815 17.6 0.815 17.6 1.395 19.61 1.395 19.61 0.815 19.84 0.815 19.84 3.685 19.41 3.685 19.41 3.215 19.365 3.215 17.605 3.215 17.605 3.685 17.37 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.105 4.59 3.105 3.09 3.335 3.09 3.335 4.59 4.795 4.59 7.185 4.59 7.185 3.56 7.415 3.56 7.415 4.59 8.435 4.59 8.925 4.59 8.925 3.39 9.155 3.39 9.155 4.59 9.65 4.59 10.225 4.59 13.33 4.59 13.33 4.345 13.56 4.345 13.56 4.59 15.06 4.59 15.37 4.59 15.37 3.875 15.605 3.875 15.605 4.59 16.345 4.59 16.345 3.875 16.58 3.875 16.58 4.59 18.39 4.59 18.39 3.875 18.62 3.875 18.62 4.585 19.365 4.585 20.43 4.585 20.43 3.875 20.66 3.875 20.66 4.59 21.28 4.59 21.28 5.49 19.365 5.49 15.06 5.49 10.225 5.49 9.65 5.49 8.435 5.49 4.795 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.96 0.45 20.96 1.165 20.73 1.165 20.73 0.45 18.72 0.45 18.72 1.165 18.49 1.165 18.49 0.45 16.535 0.45 16.535 0.64 13.34 0.64 13.34 1.37 13.11 1.37 13.11 0.45 8.535 0.45 8.535 1.37 8.305 1.37 8.305 0.45 3.455 0.45 3.455 1.37 3.225 1.37 3.225 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 1.685 0.245 1.685 0.245 1.315 0.475 1.315 0.475 1.455 2.035 1.455 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.125 1.26 4.575 1.26 4.575 3.73 4.125 3.73  ;
        POLYGON 2.615 2.63 3.895 2.63 3.895 4.02 4.795 4.02 4.795 4.36 3.665 4.36 3.665 2.86 2.615 2.86 2.615 3.685 2.385 3.685 2.385 1.26 2.715 1.26 2.715 1.6 2.615 1.6  ;
        POLYGON 6.165 3.09 8.435 3.09 8.435 3.9 8.205 3.9 8.205 3.32 6.395 3.32 6.395 3.9 6.165 3.9  ;
        POLYGON 5.375 2.63 9.65 2.63 9.65 2.86 5.375 2.86 5.375 3.73 5.145 3.73 5.145 1.26 5.695 1.26 5.695 1.6 5.375 1.6  ;
        POLYGON 6.69 2.06 9.75 2.06 9.75 1.26 9.98 1.26 9.98 2.2 10.225 2.2 10.225 4.03 9.995 4.03 9.995 2.43 9.765 2.43 9.765 2.29 6.69 2.29  ;
        POLYGON 6.145 1.6 9.29 1.6 9.29 0.8 11.685 0.8 11.685 3.1 11.455 3.1 11.455 1.03 10.64 1.03 10.64 2.06 10.41 2.06 10.41 1.03 9.52 1.03 9.52 1.83 6.375 1.83 6.375 2.06 6.145 2.06  ;
        POLYGON 11.99 1.26 12.265 1.26 12.265 3.56 11.99 3.56  ;
        POLYGON 10.87 1.26 11.1 1.26 11.1 3.22 11.245 3.22 11.245 3.8 14.83 3.8 14.83 2.415 15.06 2.415 15.06 4.03 10.87 4.03  ;
        POLYGON 12.67 2.76 14.35 2.76 14.35 1.955 15.53 1.955 15.53 1.315 15.76 1.315 15.76 1.955 19.365 1.955 19.365 2.185 14.58 2.185 14.58 3.215 12.67 3.215  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.72 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.965 2.315 4.01 2.315 4.01 2.545 3.77 2.545 3.77 2.71 2.965 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.3 2.33 17.21 2.33 17.21 2.89 16.3 2.89  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 2.89 14.825 2.89 14.825 2.47 15.055 2.47 15.055 3.27 14.71 3.27  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.48 1.58 2.48 1.58 3.27 0.71 3.27  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.125 0.845 19.45 0.845 19.45 3.685 19.125 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.96 1.495 3.96 1.495 4.59 2.055 4.59 3.005 4.59 3.005 3.56 3.235 3.56 3.235 4.59 4.835 4.59 7.245 4.59 7.245 4.49 7.475 4.49 7.475 4.59 10.445 4.59 10.445 4.49 10.675 4.49 10.675 4.59 12.49 4.59 14.33 4.59 14.33 4.005 14.67 4.005 14.67 4.59 16.37 4.59 16.37 4.005 16.71 4.005 16.71 4.59 18.135 4.59 18.465 4.59 18.465 3.48 18.695 3.48 18.695 4.59 18.895 4.59 20.205 4.59 20.205 3.875 20.435 3.875 20.435 4.59 20.72 4.59 20.72 5.49 18.895 5.49 18.135 5.49 12.49 5.49 4.835 5.49 2.055 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.72 -0.45 20.72 0.45 20.475 0.45 20.475 1.165 20.245 1.165 20.245 0.45 16.59 0.45 16.59 1.225 16.36 1.225 16.36 0.45 8.815 0.45 8.815 1.425 8.585 1.425 8.585 0.45 3.515 0.45 3.515 1.425 3.285 1.425 3.285 0.45 1.615 0.45 1.615 1.225 1.385 1.225 1.385 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.39 0.475 3.39 0.475 3.5 1.825 3.5 1.825 1.74 0.265 1.74 0.265 1.315 0.495 1.315 0.495 1.51 2.055 1.51 2.055 3.73 0.245 3.73  ;
        POLYGON 4.025 2.775 4.405 2.775 4.405 1.315 4.635 1.315 4.635 3.005 4.255 3.005 4.255 3.73 4.025 3.73  ;
        POLYGON 2.285 1.315 2.735 1.315 2.735 3.1 3.695 3.1 3.695 4.02 4.835 4.02 4.835 4.36 3.465 4.36 3.465 3.33 2.515 3.33 2.515 3.75 2.285 3.75  ;
        POLYGON 6.065 3.35 8.715 3.35 8.715 3.8 6.065 3.8  ;
        POLYGON 5.045 2.685 5.525 2.685 5.525 1.315 5.755 1.315 5.755 2.685 9.265 2.685 9.265 2.575 9.495 2.575 9.495 2.915 5.275 2.915 5.275 3.73 5.045 3.73  ;
        POLYGON 9.955 3.57 11.625 3.57 11.625 2.875 11.855 2.875 11.855 3.8 9.205 3.8 9.205 3.46 9.725 3.46 9.725 2.345 7.035 2.345 7.035 2.455 6.805 2.455 6.805 2.115 10.545 2.115 10.545 1.315 10.775 1.315 10.775 2.345 9.955 2.345  ;
        POLYGON 5.57 4.03 12.49 4.03 12.49 4.26 5.91 4.26 5.91 4.305 5.57 4.305  ;
        POLYGON 5.985 1.655 10.085 1.655 10.085 0.68 13.525 0.68 13.525 2.275 13.295 2.275 13.295 0.91 10.315 0.91 10.315 1.885 6.215 1.885 6.215 2.115 5.985 2.115  ;
        POLYGON 12.785 1.315 13.015 1.315 13.015 2.505 14.265 2.505 14.265 1.315 14.63 1.315 14.63 2.01 15.635 2.01 15.635 3.27 15.405 3.27 15.405 2.24 14.495 2.24 14.495 2.735 13.895 2.735 13.895 3.215 13.665 3.215 13.665 2.735 12.785 2.735  ;
        POLYGON 11.665 1.315 11.895 1.315 11.895 2.415 12.315 2.415 12.315 2.965 12.875 2.965 12.875 3.545 17.905 3.545 17.905 2.47 18.135 2.47 18.135 3.775 12.645 3.775 12.645 3.195 12.085 3.195 12.085 2.645 11.665 2.645  ;
        POLYGON 15.865 1.83 18.32 1.83 18.32 1.315 18.55 1.315 18.55 1.975 18.895 1.975 18.895 2.315 18.32 2.315 18.32 2.06 17.675 2.06 17.675 3.27 17.445 3.27 17.445 2.06 15.865 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.84 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.27 4.01 2.27 4.01 2.5 3.77 2.5 3.77 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.04 2.33 17.275 2.33 17.275 2.71 16.04 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.22 1.77 15.115 1.77 15.115 2.15 14.22 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.2 1.575 2.2 1.575 2.71 0.685 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.245 0.845 20.57 0.845 20.57 3.685 20.245 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.425 1.495 3.425 1.495 4.59 2.035 4.59 3.005 4.59 3.005 3.515 3.235 3.515 3.235 4.59 4.835 4.59 7.305 4.59 7.305 4.49 7.535 4.49 7.535 4.59 10.505 4.59 10.505 4.49 10.735 4.49 10.735 4.59 12.55 4.59 14.39 4.59 14.39 3.95 14.73 3.95 14.73 4.59 16.43 4.59 16.43 3.95 16.77 3.95 16.77 4.59 18.195 4.59 18.525 4.59 18.525 3.425 18.755 3.425 18.755 4.59 19.245 4.59 19.245 3.875 19.475 3.875 19.475 4.59 19.795 4.59 21.285 4.59 21.285 3.875 21.515 3.875 21.515 4.59 21.84 4.59 21.84 5.49 19.795 5.49 18.195 5.49 12.55 5.49 4.835 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.84 -0.45 21.84 0.45 21.595 0.45 21.595 1.165 21.365 1.165 21.365 0.45 19.355 0.45 19.355 1.165 19.125 1.165 19.125 0.45 16.635 0.45 16.635 1.225 16.405 1.225 16.405 0.45 8.875 0.45 8.875 1.425 8.645 1.425 8.645 0.45 3.515 0.45 3.515 1.425 3.285 1.425 3.285 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.17 0.475 3.17 0.475 3.75 0.245 3.75  ;
        POLYGON 4.025 2.73 4.405 2.73 4.405 1.315 4.635 1.315 4.635 2.96 4.255 2.96 4.255 3.685 4.025 3.685  ;
        POLYGON 2.285 1.315 2.715 1.315 2.715 3.055 3.695 3.055 3.695 3.975 4.835 3.975 4.835 4.315 3.465 4.315 3.465 3.285 2.515 3.285 2.515 3.685 2.285 3.685  ;
        POLYGON 6.065 3.35 8.775 3.35 8.775 3.8 6.065 3.8  ;
        POLYGON 5.045 2.875 5.525 2.875 5.525 1.315 5.755 1.315 5.755 2.875 9.325 2.875 9.325 2.575 9.555 2.575 9.555 3.105 5.275 3.105 5.275 3.685 5.045 3.685  ;
        POLYGON 9.265 3.46 10.605 3.46 10.605 2.345 7.035 2.345 7.035 2.455 6.805 2.455 6.805 2.115 10.605 2.115 10.605 1.315 10.835 1.315 10.835 3.57 11.685 3.57 11.685 2.875 11.915 2.875 11.915 3.8 9.265 3.8  ;
        POLYGON 5.57 4.03 12.55 4.03 12.55 4.26 5.57 4.26  ;
        POLYGON 5.985 1.655 10.145 1.655 10.145 0.68 13.79 0.68 13.79 0.91 10.375 0.91 10.375 1.885 6.215 1.885 6.215 2.115 5.985 2.115  ;
        POLYGON 12.845 1.2 15.68 1.2 15.68 2.875 15.695 2.875 15.695 3.215 15.45 3.215 15.45 1.54 13.955 1.54 13.955 3.215 13.725 3.215 13.725 1.65 12.845 1.65  ;
        POLYGON 11.725 1.315 11.955 1.315 11.955 1.88 12.935 1.88 12.935 3.455 17.965 3.455 17.965 2.415 18.195 2.415 18.195 3.685 12.705 3.685 12.705 2.11 11.725 2.11  ;
        POLYGON 15.91 1.87 18.365 1.87 18.365 1.315 18.595 1.315 18.595 1.775 19.795 1.775 19.795 2.115 17.735 2.115 17.735 3.215 17.505 3.215 17.505 2.1 15.91 2.1  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.08 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.27 4.01 2.27 4.01 2.5 3.77 2.5 3.77 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.185 2.33 17.275 2.33 17.275 2.71 16.185 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.26 1.77 15.115 1.77 15.115 2.15 14.26 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.2 1.575 2.2 1.575 2.71 0.685 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.205 2.875 22.07 2.875 22.3 2.875 22.3 1.655 20.205 1.655 20.205 0.845 20.435 0.845 20.435 1.395 22.445 1.395 22.445 0.845 22.885 0.845 22.885 3.685 22.305 3.685 22.305 3.105 22.07 3.105 20.495 3.105 20.495 3.685 20.205 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.425 1.495 3.425 1.495 4.59 2.035 4.59 3.005 4.59 3.005 3.515 3.235 3.515 3.235 4.59 4.835 4.59 7.305 4.59 7.305 4.49 7.535 4.49 7.535 4.59 10.505 4.59 10.505 4.49 10.735 4.49 10.735 4.59 12.55 4.59 14.39 4.59 14.39 3.95 14.73 3.95 14.73 4.59 16.43 4.59 16.43 3.95 16.77 3.95 16.77 4.59 18.195 4.59 18.525 4.59 18.525 3.425 18.755 3.425 18.755 4.59 19.245 4.59 19.245 3.875 19.475 3.875 19.475 4.59 21.285 4.59 21.285 3.875 21.515 3.875 21.515 4.59 22.07 4.59 23.325 4.59 23.325 3.875 23.555 3.875 23.555 4.59 24.08 4.59 24.08 5.49 22.07 5.49 18.195 5.49 12.55 5.49 4.835 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 24.08 -0.45 24.08 0.45 23.795 0.45 23.795 1.165 23.565 1.165 23.565 0.45 21.555 0.45 21.555 1.165 21.325 1.165 21.325 0.45 19.315 0.45 19.315 1.165 19.085 1.165 19.085 0.45 16.635 0.45 16.635 1.225 16.405 1.225 16.405 0.45 8.875 0.45 8.875 1.425 8.645 1.425 8.645 0.45 3.515 0.45 3.515 1.425 3.285 1.425 3.285 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.17 0.475 3.17 0.475 3.75 0.245 3.75  ;
        POLYGON 4.025 2.73 4.405 2.73 4.405 1.315 4.635 1.315 4.635 2.96 4.255 2.96 4.255 3.685 4.025 3.685  ;
        POLYGON 2.285 1.315 2.715 1.315 2.715 3.055 3.695 3.055 3.695 3.975 4.835 3.975 4.835 4.315 3.465 4.315 3.465 3.285 2.515 3.285 2.515 3.685 2.285 3.685  ;
        POLYGON 6.065 3.35 8.775 3.35 8.775 3.8 6.065 3.8  ;
        POLYGON 5.045 2.875 5.525 2.875 5.525 1.315 5.755 1.315 5.755 2.875 9.325 2.875 9.325 2.575 9.555 2.575 9.555 3.105 5.275 3.105 5.275 3.685 5.045 3.685  ;
        POLYGON 9.265 3.46 10.605 3.46 10.605 2.345 7.035 2.345 7.035 2.455 6.805 2.455 6.805 2.115 10.605 2.115 10.605 1.315 10.835 1.315 10.835 3.57 11.685 3.57 11.685 2.875 11.915 2.875 11.915 3.8 9.265 3.8  ;
        POLYGON 5.57 4.03 12.55 4.03 12.55 4.26 5.57 4.26  ;
        POLYGON 5.985 1.655 10.145 1.655 10.145 0.68 13.79 0.68 13.79 0.91 10.375 0.91 10.375 1.885 6.215 1.885 6.215 2.115 5.985 2.115  ;
        POLYGON 12.845 1.2 15.68 1.2 15.68 2.875 15.695 2.875 15.695 3.215 15.45 3.215 15.45 1.54 13.955 1.54 13.955 3.215 13.725 3.215 13.725 1.65 12.845 1.65  ;
        POLYGON 11.725 1.315 11.955 1.315 11.955 1.88 12.935 1.88 12.935 3.455 17.965 3.455 17.965 2.415 18.195 2.415 18.195 3.685 12.705 3.685 12.705 2.11 11.725 2.11  ;
        POLYGON 15.91 1.87 18.365 1.87 18.365 1.315 18.595 1.315 18.595 1.865 19.755 1.865 19.755 1.975 22.07 1.975 22.07 2.315 19.52 2.315 19.52 2.115 17.735 2.115 17.735 3.215 17.505 3.215 17.505 2.1 15.91 2.1  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.16 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 4.03 1.77 4.03 2.15 2.95 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.97 1.83 14.655 1.83 14.655 2.17 12.97 2.17  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.33 1.53 2.33 1.53 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.19 0.845 19.45 0.845 19.45 3.685 19.19 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.145 3.535 3.145 3.535 4.59 5.15 4.59 7.525 4.59 7.525 3.96 7.755 3.96 7.755 4.59 10.005 4.59 10.005 4.005 10.235 4.005 10.235 4.59 11.575 4.59 13.985 4.59 13.985 3.145 14.215 3.145 14.215 4.59 15.235 4.59 16.025 4.59 16.025 3.615 16.255 3.615 16.255 4.59 18.185 4.59 18.185 3.875 18.415 3.875 18.415 4.59 18.855 4.59 20.16 4.59 20.16 5.49 18.855 5.49 15.235 5.49 11.575 5.49 5.15 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.16 -0.45 20.16 0.45 18.315 0.45 18.315 1.165 18.085 1.165 18.085 0.45 16.475 0.45 16.475 1.265 16.245 1.265 16.245 0.45 7.635 0.45 7.635 1.245 7.405 1.245 7.405 0.45 3.435 0.45 3.435 1.245 3.205 1.245 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.325 1.135 4.555 1.135 4.555 3.785 4.325 3.785  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 2.685 3.995 2.685 3.995 4.13 5.15 4.13 5.15 4.36 3.765 4.36 3.765 2.915 2.615 2.915 2.615 3.685 2.385 3.685  ;
        POLYGON 5.445 1.135 5.675 1.135 5.675 2.11 8.47 2.11 8.47 2.34 5.675 2.34 5.675 3.785 5.445 3.785  ;
        POLYGON 6.07 1.65 7.865 1.65 7.865 0.68 10.51 0.68 10.51 0.91 8.095 0.91 8.095 1.88 6.07 1.88  ;
        POLYGON 6.81 2.57 9.785 2.57 9.785 1.315 10.015 1.315 10.015 2.975 11.135 2.975 11.135 3.315 8.765 3.315 8.765 2.8 6.81 2.8  ;
        POLYGON 5.97 3.5 8.035 3.5 8.035 3.545 11.575 3.545 11.575 4.315 11.345 4.315 11.345 3.775 7.895 3.775 7.895 3.73 6.31 3.73 6.31 4.36 5.97 4.36  ;
        POLYGON 12.74 2.4 13.495 2.4 13.495 2.685 15.235 2.685 15.235 3.785 15.005 3.785 15.005 2.915 13.495 2.915 13.495 3.685 13.265 3.685 13.265 2.63 12.51 2.63 12.51 1.655 12.025 1.655 12.025 1.26 14.215 1.26 14.215 1.6 12.74 1.6  ;
        POLYGON 10.905 0.8 15.115 0.8 15.115 1.83 16.97 1.83 16.97 2.06 14.885 2.06 14.885 1.03 11.135 1.03 11.135 1.885 12.155 1.885 12.155 3.685 11.925 3.685 11.925 2.115 10.905 2.115  ;
        POLYGON 15.585 2.515 17.365 2.515 17.365 1.315 17.595 1.315 17.595 2.39 18.855 2.39 18.855 2.73 17.455 2.73 17.455 3.215 15.585 3.215  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.72 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.075 1.77 3.975 1.77 3.975 2.15 3.075 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.435 1.21 14.97 1.21 14.97 1.59 14.665 1.59 14.665 2.115 14.435 2.115  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.24 1.39 2.24 1.39 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.125 0.845 19.45 0.845 19.45 3.685 19.125 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.895 1.595 3.895 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.615 3.535 3.615 3.535 4.59 5.295 4.59 7.475 4.59 7.475 3.615 7.705 3.615 7.705 4.59 9.875 4.59 9.875 3.83 10.105 3.83 10.105 4.59 11.445 4.59 13.855 4.59 13.855 3.515 14.085 3.515 14.085 4.59 15.105 4.59 15.895 4.59 15.895 3.045 16.125 3.045 16.125 4.59 18.105 4.59 18.105 3.875 18.335 3.875 18.335 4.59 18.775 4.59 20.145 4.59 20.145 3.875 20.375 3.875 20.375 4.59 20.72 4.59 20.72 5.49 18.775 5.49 15.105 5.49 11.445 5.49 5.295 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.72 -0.45 20.72 0.45 20.475 0.45 20.475 1.165 20.245 1.165 20.245 0.45 18.235 0.45 18.235 1.165 18.005 1.165 18.005 0.45 16.345 0.45 16.345 1.165 16.115 1.165 16.115 0.45 7.705 0.45 7.705 1.32 7.475 1.32 7.475 0.45 3.435 0.45 3.435 1.32 3.205 1.32 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.9 0.575 2.9 0.575 3.01 1.805 3.01 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.24 0.345 3.24  ;
        POLYGON 4.325 1.21 4.555 1.21 4.555 3.785 4.325 3.785  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 2.985 3.995 2.985 3.995 4.13 5.295 4.13 5.295 4.36 3.765 4.36 3.765 3.215 2.385 3.215  ;
        POLYGON 5.445 1.21 5.675 1.21 5.675 2.185 6.64 2.185 6.64 2.11 8.42 2.11 8.42 2.34 6.81 2.34 6.81 2.415 5.82 2.415 5.82 3.785 5.445 3.785  ;
        POLYGON 6.13 1.65 7.935 1.65 7.935 0.68 10.38 0.68 10.38 0.91 8.165 0.91 8.165 1.88 6.47 1.88 6.47 1.955 6.13 1.955  ;
        POLYGON 6.98 2.57 9.655 2.57 9.655 1.315 9.885 1.315 9.885 2.57 11.005 2.57 11.005 3.215 10.775 3.215 10.775 2.8 8.805 2.8 8.805 3.315 8.575 3.315 8.575 2.8 6.98 2.8  ;
        POLYGON 6.115 3.155 8.165 3.155 8.165 3.545 9.425 3.545 9.425 3.37 10.445 3.37 10.445 3.445 11.445 3.445 11.445 4.315 11.215 4.315 11.215 3.675 10.275 3.675 10.275 3.6 9.65 3.6 9.65 3.775 7.935 3.775 7.935 3.385 6.455 3.385 6.455 4.36 6.115 4.36  ;
        POLYGON 13.365 2.985 15.105 2.985 15.105 3.795 14.875 3.795 14.875 3.215 13.135 3.215 13.135 1.655 11.895 1.655 11.895 1.21 14.165 1.21 14.165 1.55 13.365 1.55  ;
        POLYGON 10.775 0.75 15.43 0.75 15.43 1.83 16.84 1.83 16.84 2.06 15.2 2.06 15.2 0.98 11.665 0.98 11.665 1.885 12.025 1.885 12.025 3.685 11.795 3.685 11.795 2.115 11.435 2.115 11.435 0.98 11.005 0.98 11.005 1.425 10.775 1.425  ;
        POLYGON 15.455 2.29 17.215 2.29 17.215 0.845 17.465 0.845 17.465 1.775 18.775 1.775 18.775 2.115 17.445 2.115 17.445 3.685 17.135 3.685 17.135 2.63 15.455 2.63  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.33 4.03 2.33 4.03 2.71 2.945 2.71  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.53 2.22 14.515 2.22 14.515 2.71 13.53 2.71  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.24 1.57 2.24 1.57 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.11 2.875 20.92 2.875 21.59 2.875 21.59 1.655 19.405 1.655 19.405 0.845 19.64 0.845 19.64 1.395 21.59 1.395 21.59 0.845 21.88 0.845 21.88 3.685 21.15 3.685 21.15 3.105 20.92 3.105 19.34 3.105 19.34 3.685 19.11 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.09 4.59 3.305 4.59 3.305 3.615 3.535 3.615 3.535 4.59 5.295 4.59 7.51 4.59 7.51 3.615 7.74 3.615 7.74 4.59 9.715 4.59 9.715 3.885 10.055 3.885 10.055 4.59 11.38 4.59 13.79 4.59 13.79 3.515 14.02 3.515 14.02 4.59 15.04 4.59 15.83 4.59 15.83 3.045 16.06 3.045 16.06 4.59 18.09 4.59 18.09 3.875 18.32 3.875 18.32 4.59 20.13 4.59 20.13 3.875 20.36 3.875 20.36 4.59 20.92 4.59 22.17 4.59 22.17 3.875 22.4 3.875 22.4 4.59 23.52 4.59 23.52 5.49 20.92 5.49 15.04 5.49 11.38 5.49 5.295 5.49 2.09 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 23 0.45 23 1.165 22.77 1.165 22.77 0.45 20.76 0.45 20.76 1.165 20.53 1.165 20.53 0.45 18.52 0.45 18.52 1.165 18.29 1.165 18.29 0.45 16.335 0.45 16.335 0.64 15.995 0.64 15.995 0.45 7.795 0.45 7.795 1.37 7.455 1.37 7.455 0.45 3.435 0.45 3.435 1.425 3.205 1.425 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.86 2.94 1.86 1.685 0.245 1.685 0.245 1.315 0.475 1.315 0.475 1.455 2.09 1.455 2.09 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.325 1.315 4.555 1.315 4.555 3.785 4.325 3.785  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.155 3.995 3.155 3.995 4.13 5.295 4.13 5.295 4.36 3.765 4.36 3.765 3.385 2.615 3.385 2.615 3.685 2.385 3.685  ;
        POLYGON 5.445 1.315 5.675 1.315 5.675 2.29 6.565 2.29 6.565 2.11 8.235 2.11 8.235 2.34 6.79 2.34 6.79 2.52 5.82 2.52 5.82 3.785 5.445 3.785  ;
        POLYGON 6 1.65 9.09 1.65 9.09 0.68 10.315 0.68 10.315 0.91 9.32 0.91 9.32 1.88 6.34 1.88 6.34 2.06 6 2.06  ;
        POLYGON 7.015 2.57 9.55 2.57 9.55 1.315 9.78 1.315 9.78 2.57 10.995 2.57 10.995 3.16 10.655 3.16 10.655 2.8 8.815 2.8 8.815 3.26 8.475 3.26 8.475 2.8 7.015 2.8  ;
        POLYGON 6.115 3.155 8.2 3.155 8.2 3.49 9.32 3.49 9.32 3.425 11.38 3.425 11.38 4.315 11.15 4.315 11.15 3.655 9.545 3.655 9.545 3.72 7.97 3.72 7.97 3.385 6.455 3.385 6.455 4.36 6.115 4.36  ;
        POLYGON 13.3 2.985 14.81 2.985 14.81 2.875 15.04 2.875 15.04 3.685 14.81 3.685 14.81 3.215 13.07 3.215 13.07 1.655 11.83 1.655 11.83 1.315 14.1 1.315 14.1 1.655 13.3 1.655  ;
        POLYGON 10.71 0.855 15.91 0.855 15.91 1.83 16.775 1.83 16.775 2.06 15.68 2.06 15.68 1.085 11.6 1.085 11.6 1.885 11.96 1.885 11.96 3.685 11.73 3.685 11.73 2.115 11.37 2.115 11.37 1.425 10.71 1.425  ;
        POLYGON 15.25 2.18 15.48 2.18 15.48 2.29 17.075 2.29 17.075 0.845 17.4 0.845 17.4 2.03 20.92 2.03 20.92 2.325 17.305 2.325 17.305 3.685 17.07 3.685 17.07 2.52 15.25 2.52  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.16 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.77 1.045 1.77 1.045 2.495 0.705 2.495  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 4.07 5.185 4.07 5.535 4.07 5.535 0.845 5.865 0.845 5.865 4.33 5.185 4.33 5.13 4.33  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.24 1.495 3.24 1.495 4.59 2.035 4.59 4.125 4.59 4.125 3.24 4.355 3.24 4.355 4.59 5.185 4.59 6.16 4.59 6.16 5.49 5.185 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.16 -0.45 6.16 0.45 4.745 0.45 4.745 0.695 4.515 0.695 4.515 0.45 1.595 0.45 1.595 1.62 1.365 1.62 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.28 0.475 1.28 0.475 2.725 1.805 2.725 1.805 1.74 2.035 1.74 2.035 2.955 0.475 2.955 0.475 3.58 0.245 3.58  ;
        POLYGON 2.385 1.28 2.715 1.28 2.715 1.795 3.83 1.795 3.83 2.495 2.615 2.495 2.615 3.58 2.385 3.58  ;
        POLYGON 3.105 2.78 4.06 2.78 4.06 1.745 4.055 1.745 4.055 0.91 3 0.91 3 0.68 4.285 0.68 4.285 1.695 5.185 1.695 5.185 2.585 4.29 2.585 4.29 3.01 3.335 3.01 3.335 3.58 3.105 3.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.21 0.97 1.21 0.97 2.795 0.71 2.795  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 3.035 5.975 3.035 6.205 3.035 6.205 1.99 5.485 1.99 5.485 0.845 5.715 0.845 5.715 1.76 6.435 1.76 6.435 3.265 5.975 3.265 5.615 3.265 5.615 4.33 5.13 4.33  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.485 1.495 3.485 1.495 4.59 2.035 4.59 4.13 4.59 4.13 3.485 4.36 3.485 4.36 4.59 5.975 4.59 6.505 4.59 6.505 3.485 6.735 3.485 6.735 4.59 7.28 4.59 7.28 5.49 5.975 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 6.855 0.45 6.855 1.63 6.625 1.63 6.625 0.45 4.595 0.45 4.595 0.96 4.365 0.96 4.365 0.45 1.595 0.45 1.595 1.645 1.365 1.645 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.305 0.475 1.305 0.475 3.025 1.805 3.025 1.805 1.985 2.035 1.985 2.035 3.255 0.475 3.255 0.475 3.825 0.245 3.825  ;
        POLYGON 2.385 1.305 2.715 1.305 2.715 2.04 3.835 2.04 3.835 2.795 3.55 2.795 3.55 2.27 2.615 2.27 2.615 3.825 2.385 3.825  ;
        POLYGON 3.11 3.025 4.065 3.025 4.065 1.41 2.955 1.41 2.955 0.68 3.295 0.68 3.295 1.18 4.295 1.18 4.295 2.22 5.975 2.22 5.975 2.56 4.295 2.56 4.295 3.255 3.34 3.255 3.34 3.825 3.11 3.825  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.035 1.05 2.035 1.05 2.735 0.71 2.735  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.68 2.95 7.115 2.95 7.345 2.95 7.345 2.04 5.63 2.04 5.63 0.77 5.86 0.77 5.86 1.81 7.87 1.81 7.87 0.77 8.1 0.77 8.1 2.04 7.575 2.04 7.575 2.98 8.05 2.98 8.05 4.25 7.82 4.25 7.82 3.21 7.115 3.21 5.91 3.21 5.91 4.25 5.68 4.25  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.27 4.59 1.27 3.44 1.5 3.44 1.5 4.59 2.095 4.59 4.28 4.59 4.28 3.44 4.51 3.44 4.51 4.59 6.7 4.59 6.7 3.44 6.93 3.44 6.93 4.59 7.115 4.59 8.89 4.59 8.89 3.44 9.12 3.44 9.12 4.59 9.52 4.59 9.52 5.49 7.115 5.49 2.095 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 9.22 0.45 9.22 1.58 8.99 1.58 8.99 0.45 6.98 0.45 6.98 1.58 6.75 1.58 6.75 0.45 4.56 0.45 4.56 1.11 4.33 1.11 4.33 0.45 1.6 0.45 1.6 1.11 1.37 1.11 1.37 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 0.77 0.48 0.77 0.48 2.965 1.755 2.965 1.755 2.035 2.095 2.035 2.095 3.195 0.48 3.195 0.48 3.78 0.25 3.78  ;
        POLYGON 2.39 2.505 3.7 2.505 3.7 2.03 2.49 2.03 2.49 0.77 2.72 0.77 2.72 1.8 3.985 1.8 3.985 2.735 2.62 2.735 2.62 3.78 2.39 3.78  ;
        POLYGON 3.26 2.98 4.215 2.98 4.215 1.57 3.21 1.57 3.21 0.77 3.44 0.77 3.44 1.34 4.445 1.34 4.445 2.27 7.115 2.27 7.115 2.5 4.445 2.5 4.445 3.21 3.49 3.21 3.49 3.78 3.26 3.78  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.77 0.99 1.77 0.99 2.56 0.65 2.56  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 2.89 6.24 2.89 6.635 2.89 6.635 0.68 6.865 0.68 6.865 4.34 6.535 4.34 6.535 3.27 6.24 3.27 5.19 3.27  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 4.02 1.495 4.02 1.495 4.59 4.385 4.59 4.735 4.59 4.735 4.04 4.965 4.04 4.965 4.59 6.24 4.59 7.28 4.59 7.28 5.49 6.24 5.49 4.385 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 5.065 0.45 5.065 0.695 4.835 0.695 4.835 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.79 1.94 2.79 1.94 1.86 2.28 1.86 2.28 3.02 0.475 3.02 0.475 4.36 0.19 4.36 0.19 0.68 0.53 0.68 0.53 0.91 0.42 0.91  ;
        POLYGON 1.555 3.3 2.51 3.3 2.51 1.63 1.5 1.63 1.5 1.4 4.385 1.4 4.385 2.615 4.155 2.615 4.155 1.63 2.74 1.63 2.74 3.64 1.555 3.64  ;
        POLYGON 4.73 1.075 5.065 1.075 5.065 1.86 6.24 1.86 6.24 2.56 5.9 2.56 5.9 2.09 4.96 2.09 4.96 3.32 4.965 3.32 4.965 3.66 4.73 3.66  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.4 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.77 0.99 1.77 0.99 2.56 0.65 2.56  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9125 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.89 6.38 2.89 6.635 2.89 6.635 0.68 6.865 0.68 6.865 4.36 6.635 4.36 6.635 3.27 6.38 3.27 6.31 3.27  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.915 1.495 3.915 1.495 4.59 4.385 4.59 4.735 4.59 4.735 3.915 4.965 3.915 4.965 4.59 6.38 4.59 7.705 4.59 7.705 3.88 7.935 3.88 7.935 4.59 8.4 4.59 8.4 5.49 6.38 5.49 4.385 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.4 -0.45 8.4 0.45 7.985 0.45 7.985 1.435 7.755 1.435 7.755 0.45 5.065 0.45 5.065 0.695 4.835 0.695 4.835 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.79 1.94 2.79 1.94 1.86 2.28 1.86 2.28 3.02 0.475 3.02 0.475 4.255 0.19 4.255 0.19 0.68 0.53 0.68 0.53 0.91 0.42 0.91  ;
        POLYGON 1.5 3.25 2.51 3.25 2.51 1.63 1.5 1.63 1.5 1.4 2.74 1.4 2.74 1.805 4.385 1.805 4.385 2.615 4.155 2.615 4.155 2.035 2.74 2.035 2.74 3.48 1.5 3.48  ;
        POLYGON 4.735 1.075 5.065 1.075 5.065 2.095 6.38 2.095 6.38 2.325 4.965 2.325 4.965 3.535 4.735 3.535  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.64 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.9 0.97 1.9 0.97 2.71 0.71 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.825 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.74 3.42 8.175 3.42 8.93 3.42 8.93 1.59 6.69 1.59 6.69 0.68 6.92 0.68 6.92 1.21 8.93 1.21 8.93 0.68 9.16 0.68 9.16 4.36 8.93 4.36 8.93 3.65 8.175 3.65 6.97 3.65 6.97 4.36 6.74 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.32 4.59 1.32 4.06 1.55 4.06 1.55 4.59 4.44 4.59 4.79 4.59 4.79 4.06 5.02 4.06 5.02 4.59 7.76 4.59 7.76 3.88 7.99 3.88 7.99 4.59 8.175 4.59 9.95 4.59 9.95 3.88 10.18 3.88 10.18 4.59 10.64 4.59 10.64 5.49 8.175 5.49 4.44 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.64 -0.45 10.64 0.45 10.28 0.45 10.28 1.435 10.05 1.435 10.05 0.45 8.04 0.45 8.04 0.965 7.81 0.965 7.81 0.45 5.12 0.45 5.12 0.695 4.89 0.695 4.89 0.45 1.65 0.45 1.65 0.965 1.42 0.965 1.42 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.94 1.275 2.94 1.275 2.425 2.05 2.425 2.05 1.9 2.335 1.9 2.335 2.655 1.505 2.655 1.505 3.17 0.585 3.17 0.585 4.345 0.245 4.345 0.245 0.68 0.585 0.68 0.585 0.91 0.475 0.91  ;
        POLYGON 1.555 3.395 2.565 3.395 2.565 1.63 1.555 1.63 1.555 1.4 4.44 1.4 4.44 2.71 4.21 2.71 4.21 1.63 2.795 1.63 2.795 3.625 1.555 3.625  ;
        POLYGON 4.79 1.075 5.12 1.075 5.12 2.19 8.175 2.19 8.175 2.42 5.02 2.42 5.02 3.68 4.79 3.68  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.2 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.77 0.97 1.77 0.97 2.56 0.63 2.56  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.23 2.89 10.295 2.89 10.69 2.89 10.69 0.68 10.92 0.68 10.92 4.36 10.59 4.36 10.59 3.27 10.295 3.27 10.23 3.27  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.84 4.59 4.44 4.59 8.44 4.59 10.295 4.59 11.2 4.59 11.2 5.49 10.295 5.49 8.44 5.49 4.44 5.49 0 5.49 0 4.59 1.61 4.59 1.61 3.88 4.44 3.88 8.44 3.88 9.02 3.88 9.02 4.22 8.44 4.22 4.44 4.22 1.84 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.2 -0.45 11.2 0.45 9.12 0.45 9.12 0.695 8.89 0.695 8.89 0.45 5.12 0.45 5.12 0.69 4.89 0.69 4.89 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.4 2.79 1.2 2.79 1.2 2.33 1.995 2.33 1.995 1.86 2.335 1.86 2.335 2.56 1.43 2.56 1.43 3.02 0.475 3.02 0.475 4.22 0.17 4.22 0.17 0.68 0.53 0.68 0.53 0.91 0.4 0.91  ;
        POLYGON 1.555 3.215 4.21 3.215 4.21 1.63 1.555 1.63 1.555 1.4 4.44 1.4 4.44 3.445 1.555 3.445  ;
        POLYGON 4.79 1.07 5.12 1.07 5.12 1.86 6.335 1.86 6.335 2.56 5.995 2.56 5.995 2.09 5.02 2.09 5.02 3.5 4.79 3.5  ;
        POLYGON 5.61 2.79 6.565 2.79 6.565 1.63 5.61 1.63 5.61 1.07 5.84 1.07 5.84 1.4 8.44 1.4 8.44 2.615 8.21 2.615 8.21 1.63 6.795 1.63 6.795 3.02 5.84 3.02 5.84 3.5 5.61 3.5  ;
        POLYGON 8.79 1.075 9.12 1.075 9.12 1.86 10.295 1.86 10.295 2.56 9.955 2.56 9.955 2.09 9.02 2.09 9.02 3.5 8.79 3.5  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.77 0.99 1.77 0.99 2.56 0.65 2.56  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9125 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.23 1.21 10.635 1.21 10.635 0.68 10.865 0.68 10.865 4.36 10.635 4.36 10.635 1.59 10.23 1.59  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.915 1.495 3.915 1.495 4.59 4.385 4.59 4.735 4.59 4.735 3.915 4.965 3.915 4.965 4.59 8.385 4.59 8.735 4.59 8.735 3.915 8.965 3.915 8.965 4.59 10.38 4.59 11.705 4.59 11.705 3.88 11.935 3.88 11.935 4.59 12.32 4.59 12.32 5.49 10.38 5.49 8.385 5.49 4.385 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 11.985 0.45 11.985 1.435 11.755 1.435 11.755 0.45 9.065 0.45 9.065 0.695 8.835 0.695 8.835 0.45 5.065 0.45 5.065 0.69 4.835 0.69 4.835 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.79 1.94 2.79 1.94 1.86 2.28 1.86 2.28 3.02 0.475 3.02 0.475 4.255 0.19 4.255 0.19 0.68 0.53 0.68 0.53 0.91 0.42 0.91  ;
        POLYGON 1.5 3.25 2.51 3.25 2.51 1.63 1.5 1.63 1.5 1.4 4.385 1.4 4.385 2.615 4.155 2.615 4.155 1.63 2.74 1.63 2.74 3.48 1.5 3.48  ;
        POLYGON 4.735 1.07 5.065 1.07 5.065 1.86 6.28 1.86 6.28 2.56 5.94 2.56 5.94 2.09 4.965 2.09 4.965 3.535 4.735 3.535  ;
        POLYGON 5.555 2.79 6.51 2.79 6.51 1.63 5.555 1.63 5.555 1.07 5.785 1.07 5.785 1.4 8.385 1.4 8.385 2.615 8.155 2.615 8.155 1.63 6.74 1.63 6.74 3.02 5.785 3.02 5.785 3.535 5.555 3.535  ;
        POLYGON 8.735 1.075 9.065 1.075 9.065 2.095 10.38 2.095 10.38 2.325 8.965 2.325 8.965 3.535 8.735 3.535  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.14 0.99 1.14 0.99 1.84 0.65 1.84  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.565 2.875 11.995 2.875 12.225 2.875 12.225 1.655 10.565 1.655 10.565 0.845 10.795 0.845 10.795 1.425 12.47 1.425 12.47 0.845 13.035 0.845 13.035 1.655 12.455 1.655 12.455 2.875 12.935 2.875 12.935 3.685 12.705 3.685 12.705 3.105 11.995 3.105 10.795 3.105 10.795 3.685 10.565 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.71 1.495 3.71 1.495 4.59 4.315 4.59 4.665 4.59 4.665 3.71 4.895 3.71 4.895 4.59 8.315 4.59 8.665 4.59 8.665 3.71 8.895 3.71 8.895 4.59 11.585 4.59 11.585 3.875 11.815 3.875 11.815 4.59 11.995 4.59 13.825 4.59 13.825 3.875 14.055 3.875 14.055 4.59 14.56 4.59 14.56 5.49 11.995 5.49 8.315 5.49 4.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 14.155 0.45 14.155 1.165 13.925 1.165 13.925 0.45 11.915 0.45 11.915 1.165 11.685 1.165 11.685 0.45 8.995 0.45 8.995 0.935 8.765 0.935 8.765 0.45 4.995 0.45 4.995 0.935 4.765 0.935 4.765 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.53 1.87 2.53 1.87 2.06 2.21 2.06 2.21 2.76 0.475 2.76 0.475 4.05 0.19 4.05 0.19 0.68 0.53 0.68 0.53 0.91 0.42 0.91  ;
        POLYGON 1.485 2.99 4.085 2.99 4.085 1.715 1.43 1.715 1.43 1.485 4.315 1.485 4.315 3.33 1.485 3.33  ;
        POLYGON 4.665 1.315 4.995 1.315 4.995 1.83 6.21 1.83 6.21 2.53 5.87 2.53 5.87 2.06 4.895 2.06 4.895 3.33 4.665 3.33  ;
        POLYGON 5.485 2.76 8.085 2.76 8.085 1.6 5.43 1.6 5.43 1.37 8.315 1.37 8.315 2.99 5.715 2.99 5.715 3.33 5.485 3.33  ;
        POLYGON 8.665 1.315 8.995 1.315 8.995 1.975 11.995 1.975 11.995 2.315 8.895 2.315 8.895 3.33 8.665 3.33  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.12 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.58 0.71 2.58  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.545 0.84 14.97 0.84 14.97 4.36 14.545 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.27 4.59 1.27 3.895 1.5 3.895 1.5 4.59 4.39 4.59 4.74 4.59 4.74 3.895 4.97 3.895 4.97 4.59 8.39 4.59 8.74 4.59 8.74 3.895 8.97 3.895 8.97 4.59 12.395 4.59 12.745 4.59 12.745 3.895 12.975 3.895 12.975 4.59 14.195 4.59 15.12 4.59 15.12 5.49 14.195 5.49 12.395 5.49 8.39 5.49 4.39 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.12 -0.45 15.12 0.45 13.075 0.45 13.075 0.69 12.845 0.69 12.845 0.45 9.07 0.45 9.07 0.93 8.84 0.93 8.84 0.45 5.07 0.45 5.07 0.93 4.84 0.93 4.84 0.45 1.6 0.45 1.6 0.965 1.37 0.965 1.37 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.425 2.81 1.245 2.81 1.245 2.77 2 2.77 2 2.19 2.23 2.19 2.23 3 1.375 3 1.375 3.04 0.48 3.04 0.48 4.235 0.195 4.235 0.195 0.68 0.535 0.68 0.535 0.91 0.425 0.91  ;
        POLYGON 1.505 3.23 2.46 3.23 2.46 1.63 1.505 1.63 1.505 1.4 4.39 1.4 4.39 2.58 4.16 2.58 4.16 1.63 2.69 1.63 2.69 3.46 1.505 3.46  ;
        POLYGON 4.74 1.31 5.07 1.31 5.07 2.35 6 2.35 6 1.77 6.23 1.77 6.23 2.58 4.97 2.58 4.97 3.515 4.74 3.515  ;
        POLYGON 5.56 2.81 6.46 2.81 6.46 1.54 5.845 1.54 5.845 1.595 5.505 1.595 5.505 1.31 8.39 1.31 8.39 2.58 8.16 2.58 8.16 1.54 6.69 1.54 6.69 3.04 5.79 3.04 5.79 3.515 5.56 3.515  ;
        POLYGON 8.74 1.31 9.07 1.31 9.07 2.35 10 2.35 10 1.77 10.23 1.77 10.23 2.58 8.97 2.58 8.97 3.515 8.74 3.515  ;
        POLYGON 9.56 2.81 10.46 2.81 10.46 1.54 9.845 1.54 9.845 1.595 9.505 1.595 9.505 1.31 12.395 1.31 12.395 2.58 12.165 2.58 12.165 1.54 10.69 1.54 10.69 3.04 9.79 3.04 9.79 3.515 9.56 3.515  ;
        POLYGON 12.745 1.07 13.075 1.07 13.075 1.77 14.195 1.77 14.195 2.58 13.965 2.58 13.965 2 12.975 2 12.975 3.515 12.745 3.515  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 16.24 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.77 0.99 1.77 0.99 2.57 0.65 2.57  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.53 4.07 14.535 4.07 14.535 3.135 15.125 3.135 15.355 3.135 15.355 1.82 14.635 1.82 14.635 0.845 14.865 0.845 14.865 1.59 15.585 1.59 15.585 3.365 15.125 3.365 14.765 3.365 14.765 4.36 13.53 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.925 1.495 3.925 1.495 4.59 4.385 4.59 4.735 4.59 4.735 3.925 4.965 3.925 4.965 4.59 8.385 4.59 8.735 4.59 8.735 3.925 8.965 3.925 8.965 4.59 12.385 4.59 12.735 4.59 12.735 3.925 12.965 3.925 12.965 4.59 15.125 4.59 15.655 4.59 15.655 3.585 15.885 3.585 15.885 4.59 16.24 4.59 16.24 5.49 15.125 5.49 12.385 5.49 8.385 5.49 4.385 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 16.24 -0.45 16.24 0.45 15.985 0.45 15.985 1.435 15.755 1.435 15.755 0.45 13.065 0.45 13.065 0.695 12.835 0.695 12.835 0.45 9.065 0.45 9.065 0.92 8.835 0.92 8.835 0.45 5.065 0.45 5.065 0.69 4.835 0.69 4.835 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.8 1.995 2.8 1.995 2.22 2.225 2.22 2.225 3.03 0.475 3.03 0.475 4.265 0.19 4.265 0.19 0.68 0.53 0.68 0.53 0.91 0.42 0.91  ;
        POLYGON 1.5 3.26 4.155 3.26 4.155 1.63 1.5 1.63 1.5 1.4 4.385 1.4 4.385 3.49 1.5 3.49  ;
        POLYGON 4.735 1.07 5.065 1.07 5.065 1.815 6.225 1.815 6.225 2.625 4.965 2.625 4.965 3.545 4.735 3.545  ;
        POLYGON 5.555 2.855 8.155 2.855 8.155 1.585 5.555 1.585 5.555 1.07 5.785 1.07 5.785 1.355 8.385 1.355 8.385 3.085 5.785 3.085 5.785 3.545 5.555 3.545  ;
        POLYGON 8.735 1.3 9.065 1.3 9.065 1.815 10.225 1.815 10.225 2.625 8.965 2.625 8.965 3.545 8.735 3.545  ;
        POLYGON 9.555 2.855 12.155 2.855 12.155 1.585 9.5 1.585 9.5 1.355 12.385 1.355 12.385 3.085 9.785 3.085 9.785 3.545 9.555 3.545  ;
        POLYGON 12.735 1.075 13.065 1.075 13.065 2.05 15.125 2.05 15.125 2.39 12.965 2.39 12.965 3.545 12.735 3.545  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 18.48 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.77 1 1.77 1 2.595 0.66 2.595  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.825 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.695 2.89 16.13 2.89 16.36 2.89 16.36 1.9 14.645 1.9 14.645 0.68 14.875 0.68 14.875 1.67 16.885 1.67 16.885 0.68 17.115 0.68 17.115 1.9 16.59 1.9 16.59 2.89 16.965 2.89 16.965 4.36 16.735 4.36 16.735 3.12 16.13 3.12 14.97 3.12 14.97 4.36 14.695 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.275 4.59 1.275 3.93 1.505 3.93 1.505 4.59 4.395 4.59 4.745 4.59 4.745 3.93 4.975 3.93 4.975 4.59 8.395 4.59 8.745 4.59 8.745 3.93 8.975 3.93 8.975 4.59 12.395 4.59 12.745 4.59 12.745 3.93 12.975 3.93 12.975 4.59 15.715 4.59 15.715 3.88 15.945 3.88 15.945 4.59 16.13 4.59 17.905 4.59 17.905 3.88 18.135 3.88 18.135 4.59 18.48 4.59 18.48 5.49 16.13 5.49 12.395 5.49 8.395 5.49 4.395 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 18.48 -0.45 18.48 0.45 18.235 0.45 18.235 1.44 18.005 1.44 18.005 0.45 15.995 0.45 15.995 1.44 15.765 1.44 15.765 0.45 13.075 0.45 13.075 0.695 12.845 0.695 12.845 0.45 9.075 0.45 9.075 0.965 8.845 0.965 8.845 0.45 5.075 0.45 5.075 0.97 4.845 0.97 4.845 0.45 1.605 0.45 1.605 0.97 1.375 0.97 1.375 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.43 2.825 1.32 2.825 1.32 2.805 1.95 2.805 1.95 1.895 2.29 1.895 2.29 3.035 1.415 3.035 1.415 3.055 0.485 3.055 0.485 4.27 0.2 4.27 0.2 0.685 0.54 0.685 0.54 0.915 0.43 0.915  ;
        POLYGON 1.51 3.265 2.52 3.265 2.52 1.635 1.51 1.635 1.51 1.405 4.395 1.405 4.395 2.65 4.165 2.65 4.165 1.635 2.75 1.635 2.75 3.495 1.51 3.495  ;
        POLYGON 4.745 1.35 5.075 1.35 5.075 1.895 6.29 1.895 6.29 2.595 5.95 2.595 5.95 2.125 4.975 2.125 4.975 3.55 4.745 3.55  ;
        POLYGON 5.565 2.825 6.52 2.825 6.52 1.635 5.51 1.635 5.51 1.405 8.395 1.405 8.395 2.65 8.165 2.65 8.165 1.635 6.75 1.635 6.75 3.055 5.795 3.055 5.795 3.55 5.565 3.55  ;
        POLYGON 8.745 1.345 9.075 1.345 9.075 1.895 10.29 1.895 10.29 2.595 9.95 2.595 9.95 2.125 8.975 2.125 8.975 3.55 8.745 3.55  ;
        POLYGON 9.565 2.825 10.52 2.825 10.52 1.63 9.51 1.63 9.51 1.4 10.75 1.4 10.75 1.84 12.395 1.84 12.395 2.65 12.165 2.65 12.165 2.07 10.75 2.07 10.75 3.055 9.795 3.055 9.795 3.55 9.565 3.55  ;
        POLYGON 12.745 1.075 13.075 1.075 13.075 2.13 16.13 2.13 16.13 2.36 12.975 2.36 12.975 3.55 12.745 3.55  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__endcap
  CLASS gf180mcu_fd_sc_mcu9t5v0__endcap PRE ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__endcap 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 1.12 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.23 4.59 0.23 2.34 0.85 2.34 0.85 4.59 1.12 4.59 1.12 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 1.12 -0.45 1.12 0.45 0.85 0.45 0.85 1.53 0.23 1.53 0.23 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__endcap
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_1
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 0.56 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.56 4.59 0.56 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 0.56 -0.45 0.56 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_2
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 1.12 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.12 4.59 1.12 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 1.12 -0.45 1.12 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.24 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.24 4.59 2.24 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.24 -0.45 2.24 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 4.48 4.59 4.48 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_8
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 8.96 4.59 8.96 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_16
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 17.92 4.59 17.92 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_32
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_64 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 35.84 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 35.84 4.59 35.84 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 35.84 -0.45 35.84 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_64
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.24 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.97 4.59 1.765 4.59 1.765 3.55 1.995 3.55 1.995 4.59 2.24 4.59 2.24 5.49 1.995 5.49 0.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.24 -0.45 2.24 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.83 0.97 1.83 0.97 2.06 0.475 2.06 0.475 4.36 0.245 4.36  ;
        POLYGON 1.27 2.47 1.765 2.47 1.765 0.68 1.995 0.68 1.995 2.7 1.27 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.97 4.59 1.765 4.59 1.765 3.55 1.995 3.55 1.995 4.59 3.21 4.59 4.005 4.59 4.005 3.55 4.235 3.55 4.235 4.59 4.48 4.59 4.48 5.49 4.235 5.49 3.21 5.49 1.995 5.49 0.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.83 0.97 1.83 0.97 2.06 0.475 2.06 0.475 4.36 0.245 4.36  ;
        POLYGON 1.27 2.47 1.765 2.47 1.765 0.68 1.995 0.68 1.995 2.7 1.27 2.7  ;
        POLYGON 2.485 1.83 3.21 1.83 3.21 2.06 2.715 2.06 2.715 4.36 2.485 4.36  ;
        POLYGON 3.51 2.47 4.005 2.47 4.005 0.68 4.235 0.68 4.235 2.7 3.51 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_8
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.97 4.59 1.765 4.59 1.765 3.55 1.995 3.55 1.995 4.59 3.21 4.59 4.005 4.59 4.005 3.55 4.235 3.55 4.235 4.59 5.45 4.59 6.245 4.59 6.245 3.55 6.475 3.55 6.475 4.59 7.69 4.59 8.485 4.59 8.485 3.55 8.715 3.55 8.715 4.59 8.96 4.59 8.96 5.49 8.715 5.49 7.69 5.49 6.475 5.49 5.45 5.49 4.235 5.49 3.21 5.49 1.995 5.49 0.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.83 0.97 1.83 0.97 2.06 0.475 2.06 0.475 4.36 0.245 4.36  ;
        POLYGON 1.27 2.47 1.765 2.47 1.765 0.68 1.995 0.68 1.995 2.7 1.27 2.7  ;
        POLYGON 2.485 1.83 3.21 1.83 3.21 2.06 2.715 2.06 2.715 4.36 2.485 4.36  ;
        POLYGON 3.51 2.47 4.005 2.47 4.005 0.68 4.235 0.68 4.235 2.7 3.51 2.7  ;
        POLYGON 4.725 1.83 5.45 1.83 5.45 2.06 4.955 2.06 4.955 4.36 4.725 4.36  ;
        POLYGON 5.75 2.47 6.245 2.47 6.245 0.68 6.475 0.68 6.475 2.7 5.75 2.7  ;
        POLYGON 6.965 1.83 7.69 1.83 7.69 2.06 7.195 2.06 7.195 4.36 6.965 4.36  ;
        POLYGON 7.99 2.47 8.485 2.47 8.485 0.68 8.715 0.68 8.715 2.7 7.99 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_16
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.97 4.59 1.765 4.59 1.765 3.55 1.995 3.55 1.995 4.59 3.21 4.59 4.005 4.59 4.005 3.55 4.235 3.55 4.235 4.59 5.45 4.59 6.245 4.59 6.245 3.55 6.475 3.55 6.475 4.59 7.69 4.59 8.485 4.59 8.485 3.55 8.715 3.55 8.715 4.59 9.93 4.59 10.725 4.59 10.725 3.55 10.955 3.55 10.955 4.59 12.17 4.59 12.965 4.59 12.965 3.55 13.195 3.55 13.195 4.59 14.41 4.59 15.205 4.59 15.205 3.55 15.435 3.55 15.435 4.59 16.65 4.59 17.445 4.59 17.445 3.55 17.675 3.55 17.675 4.59 17.92 4.59 17.92 5.49 17.675 5.49 16.65 5.49 15.435 5.49 14.41 5.49 13.195 5.49 12.17 5.49 10.955 5.49 9.93 5.49 8.715 5.49 7.69 5.49 6.475 5.49 5.45 5.49 4.235 5.49 3.21 5.49 1.995 5.49 0.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.83 0.97 1.83 0.97 2.06 0.475 2.06 0.475 4.36 0.245 4.36  ;
        POLYGON 1.325 1.26 1.765 1.26 1.765 0.68 1.995 0.68 1.995 1.49 1.555 1.49 1.555 2.755 1.325 2.755  ;
        POLYGON 2.485 1.83 3.21 1.83 3.21 2.06 2.715 2.06 2.715 4.36 2.485 4.36  ;
        POLYGON 3.565 1.26 4.005 1.26 4.005 0.68 4.235 0.68 4.235 1.49 3.795 1.49 3.795 2.755 3.565 2.755  ;
        POLYGON 4.725 1.83 5.45 1.83 5.45 2.06 4.955 2.06 4.955 4.36 4.725 4.36  ;
        POLYGON 5.805 1.26 6.245 1.26 6.245 0.68 6.475 0.68 6.475 1.49 6.035 1.49 6.035 2.755 5.805 2.755  ;
        POLYGON 6.965 1.83 7.69 1.83 7.69 2.06 7.195 2.06 7.195 4.36 6.965 4.36  ;
        POLYGON 8.045 1.26 8.485 1.26 8.485 0.68 8.715 0.68 8.715 1.49 8.275 1.49 8.275 2.755 8.045 2.755  ;
        POLYGON 9.205 1.83 9.93 1.83 9.93 2.06 9.435 2.06 9.435 4.36 9.205 4.36  ;
        POLYGON 10.285 1.26 10.725 1.26 10.725 0.68 10.955 0.68 10.955 1.49 10.515 1.49 10.515 2.755 10.285 2.755  ;
        POLYGON 11.445 1.83 12.17 1.83 12.17 2.06 11.675 2.06 11.675 4.36 11.445 4.36  ;
        POLYGON 12.525 1.26 12.965 1.26 12.965 0.68 13.195 0.68 13.195 1.49 12.755 1.49 12.755 2.755 12.525 2.755  ;
        POLYGON 13.685 1.83 14.41 1.83 14.41 2.06 13.915 2.06 13.915 4.36 13.685 4.36  ;
        POLYGON 14.765 1.26 15.205 1.26 15.205 0.68 15.435 0.68 15.435 1.49 14.995 1.49 14.995 2.755 14.765 2.755  ;
        POLYGON 15.925 1.83 16.65 1.83 16.65 2.06 16.155 2.06 16.155 4.36 15.925 4.36  ;
        POLYGON 17.005 1.26 17.445 1.26 17.445 0.68 17.675 0.68 17.675 1.49 17.235 1.49 17.235 2.755 17.005 2.755  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_32
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_64 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 35.84 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.97 4.59 1.765 4.59 1.765 3.55 1.995 3.55 1.995 4.59 3.21 4.59 4.005 4.59 4.005 3.55 4.235 3.55 4.235 4.59 5.45 4.59 6.245 4.59 6.245 3.55 6.475 3.55 6.475 4.59 7.69 4.59 8.485 4.59 8.485 3.55 8.715 3.55 8.715 4.59 9.93 4.59 10.725 4.59 10.725 3.55 10.955 3.55 10.955 4.59 12.17 4.59 12.965 4.59 12.965 3.55 13.195 3.55 13.195 4.59 14.41 4.59 15.205 4.59 15.205 3.55 15.435 3.55 15.435 4.59 16.65 4.59 17.445 4.59 17.445 3.55 17.675 3.55 17.675 4.59 18.89 4.59 19.685 4.59 19.685 3.55 19.915 3.55 19.915 4.59 21.13 4.59 21.925 4.59 21.925 3.55 22.155 3.55 22.155 4.59 23.37 4.59 24.165 4.59 24.165 3.55 24.395 3.55 24.395 4.59 25.61 4.59 26.405 4.59 26.405 3.55 26.635 3.55 26.635 4.59 27.85 4.59 28.645 4.59 28.645 3.55 28.875 3.55 28.875 4.59 30.09 4.59 30.885 4.59 30.885 3.55 31.115 3.55 31.115 4.59 32.33 4.59 33.125 4.59 33.125 3.55 33.355 3.55 33.355 4.59 34.57 4.59 35.365 4.59 35.365 3.55 35.595 3.55 35.595 4.59 35.84 4.59 35.84 5.49 35.595 5.49 34.57 5.49 33.355 5.49 32.33 5.49 31.115 5.49 30.09 5.49 28.875 5.49 27.85 5.49 26.635 5.49 25.61 5.49 24.395 5.49 23.37 5.49 22.155 5.49 21.13 5.49 19.915 5.49 18.89 5.49 17.675 5.49 16.65 5.49 15.435 5.49 14.41 5.49 13.195 5.49 12.17 5.49 10.955 5.49 9.93 5.49 8.715 5.49 7.69 5.49 6.475 5.49 5.45 5.49 4.235 5.49 3.21 5.49 1.995 5.49 0.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 35.84 -0.45 35.84 0.45 34.075 0.45 34.075 1.49 33.845 1.49 33.845 0.45 31.835 0.45 31.835 1.49 31.605 1.49 31.605 0.45 29.595 0.45 29.595 1.49 29.365 1.49 29.365 0.45 27.355 0.45 27.355 1.49 27.125 1.49 27.125 0.45 25.115 0.45 25.115 1.49 24.885 1.49 24.885 0.45 22.875 0.45 22.875 1.49 22.645 1.49 22.645 0.45 20.635 0.45 20.635 1.49 20.405 1.49 20.405 0.45 18.395 0.45 18.395 1.49 18.165 1.49 18.165 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.83 0.97 1.83 0.97 2.06 0.475 2.06 0.475 4.36 0.245 4.36  ;
        POLYGON 1.325 1.26 1.765 1.26 1.765 0.68 1.995 0.68 1.995 1.49 1.555 1.49 1.555 2.755 1.325 2.755  ;
        POLYGON 2.485 1.83 3.21 1.83 3.21 2.06 2.715 2.06 2.715 4.36 2.485 4.36  ;
        POLYGON 3.565 1.26 4.005 1.26 4.005 0.68 4.235 0.68 4.235 1.49 3.795 1.49 3.795 2.755 3.565 2.755  ;
        POLYGON 4.725 1.83 5.45 1.83 5.45 2.06 4.955 2.06 4.955 4.36 4.725 4.36  ;
        POLYGON 5.805 1.26 6.245 1.26 6.245 0.68 6.475 0.68 6.475 1.49 6.035 1.49 6.035 2.755 5.805 2.755  ;
        POLYGON 6.965 1.83 7.69 1.83 7.69 2.06 7.195 2.06 7.195 4.36 6.965 4.36  ;
        POLYGON 8.045 1.26 8.485 1.26 8.485 0.68 8.715 0.68 8.715 1.49 8.275 1.49 8.275 2.755 8.045 2.755  ;
        POLYGON 9.205 1.83 9.93 1.83 9.93 2.06 9.435 2.06 9.435 4.36 9.205 4.36  ;
        POLYGON 10.285 1.26 10.725 1.26 10.725 0.68 10.955 0.68 10.955 1.49 10.515 1.49 10.515 2.755 10.285 2.755  ;
        POLYGON 11.445 1.83 12.17 1.83 12.17 2.06 11.675 2.06 11.675 4.36 11.445 4.36  ;
        POLYGON 12.525 1.26 12.965 1.26 12.965 0.68 13.195 0.68 13.195 1.49 12.755 1.49 12.755 2.755 12.525 2.755  ;
        POLYGON 13.685 1.83 14.41 1.83 14.41 2.06 13.915 2.06 13.915 4.36 13.685 4.36  ;
        POLYGON 14.765 1.26 15.205 1.26 15.205 0.68 15.435 0.68 15.435 1.49 14.995 1.49 14.995 2.755 14.765 2.755  ;
        POLYGON 15.925 1.83 16.65 1.83 16.65 2.06 16.155 2.06 16.155 4.36 15.925 4.36  ;
        POLYGON 17.005 1.26 17.445 1.26 17.445 0.68 17.675 0.68 17.675 1.49 17.235 1.49 17.235 2.755 17.005 2.755  ;
        POLYGON 18.165 1.83 18.89 1.83 18.89 2.06 18.395 2.06 18.395 4.36 18.165 4.36  ;
        POLYGON 19.245 1.26 19.685 1.26 19.685 0.68 19.915 0.68 19.915 1.49 19.475 1.49 19.475 2.755 19.245 2.755  ;
        POLYGON 20.405 1.83 21.13 1.83 21.13 2.06 20.635 2.06 20.635 4.36 20.405 4.36  ;
        POLYGON 21.485 1.26 21.925 1.26 21.925 0.68 22.155 0.68 22.155 1.49 21.715 1.49 21.715 2.755 21.485 2.755  ;
        POLYGON 22.645 1.83 23.37 1.83 23.37 2.06 22.875 2.06 22.875 4.36 22.645 4.36  ;
        POLYGON 23.725 1.26 24.165 1.26 24.165 0.68 24.395 0.68 24.395 1.49 23.955 1.49 23.955 2.755 23.725 2.755  ;
        POLYGON 24.885 1.83 25.61 1.83 25.61 2.06 25.115 2.06 25.115 4.36 24.885 4.36  ;
        POLYGON 25.965 1.26 26.405 1.26 26.405 0.68 26.635 0.68 26.635 1.49 26.195 1.49 26.195 2.755 25.965 2.755  ;
        POLYGON 27.125 1.83 27.85 1.83 27.85 2.06 27.355 2.06 27.355 4.36 27.125 4.36  ;
        POLYGON 28.205 1.26 28.645 1.26 28.645 0.68 28.875 0.68 28.875 1.49 28.435 1.49 28.435 2.755 28.205 2.755  ;
        POLYGON 29.365 1.83 30.09 1.83 30.09 2.06 29.595 2.06 29.595 4.36 29.365 4.36  ;
        POLYGON 30.445 1.26 30.885 1.26 30.885 0.68 31.115 0.68 31.115 1.49 30.675 1.49 30.675 2.755 30.445 2.755  ;
        POLYGON 31.605 1.83 32.33 1.83 32.33 2.06 31.835 2.06 31.835 4.36 31.605 4.36  ;
        POLYGON 32.685 1.26 33.125 1.26 33.125 0.68 33.355 0.68 33.355 1.49 32.915 1.49 32.915 2.755 32.685 2.755  ;
        POLYGON 33.845 1.83 34.57 1.83 34.57 2.06 34.075 2.06 34.075 4.36 33.845 4.36  ;
        POLYGON 34.925 1.26 35.365 1.26 35.365 0.68 35.595 0.68 35.595 1.49 35.155 1.49 35.155 2.755 34.925 2.755  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_64
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__filltie
  CLASS core WELLTAP ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__filltie 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 1.12 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.33 4.59 0.33 2.34 0.71 2.34 0.71 4.59 1.12 4.59 1.12 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 1.12 -0.45 1.12 0.45 0.71 0.45 0.71 1.91 0.33 1.91 0.33 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__filltie
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__hold
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__hold 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN Z
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.4896 ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.415 3.95 1.415 3.95 2.575 3.51 2.575 3.51 1.645 0.575 1.645 0.575 3.605 0.245 3.605  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 3.225 4.59 3.225 3.265 3.455 3.265 3.455 4.59 4.575 4.59 5.04 4.59 5.04 5.49 4.575 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 3.455 0.45 3.455 1.185 3.225 1.185 3.225 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.51 1.875 2.85 1.875 2.85 2.805 4.345 2.805 4.345 0.845 4.575 0.845 4.575 4.075 4.245 4.075 4.245 3.035 2.51 3.035  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__hold
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 16.8 BY 5.04 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.22 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.35 1.77 11.715 1.77 11.715 2.71 11.35 2.71  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 1.77 2.09 1.77 2.09 2.265 1.21 2.265  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.915 1.77 0.915 2.265 0.41 2.265 0.41 2.71 0.15 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2452 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.83 3.39 16.245 3.39 16.245 1.59 15.83 1.59 15.83 1.21 16.245 1.21 16.245 0.795 16.475 0.795 16.475 4.2 16.195 4.2 16.195 3.83 15.83 3.83  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.675 4.59 0.675 3.39 0.905 3.39 0.905 4.59 2.715 4.59 5.805 4.59 5.805 3.39 6.035 3.39 6.035 4.59 8.335 4.59 8.665 4.59 8.665 3.39 8.895 3.39 8.895 4.59 9.39 4.59 12.245 4.59 12.245 3.39 12.475 3.39 12.475 4.59 12.915 4.59 15.175 4.59 15.175 3.39 15.405 3.39 15.405 4.59 15.74 4.59 16.8 4.59 16.8 5.49 15.74 5.49 12.915 5.49 9.39 5.49 8.335 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 16.8 -0.45 16.8 0.45 15.355 0.45 15.355 1.605 15.125 1.605 15.125 0.45 14.635 0.45 14.635 1.135 14.405 1.135 14.405 0.45 12.395 0.45 12.395 1.135 12.165 1.135 12.165 0.45 8.995 0.45 8.995 1.135 8.765 1.135 8.765 0.45 6.035 0.45 6.035 1.135 5.805 1.135 5.805 0.45 1.65 0.45 1.65 1.08 1.31 1.08 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.795 0.475 0.795 0.475 1.31 2.485 1.31 2.485 0.795 2.715 0.795 2.715 1.54 0.245 1.54  ;
        POLYGON 3.445 1.79 3.675 1.79 3.675 2.47 6.925 2.47 6.925 0.795 7.155 0.795 7.155 3.9 6.825 3.9 6.825 2.7 3.445 2.7  ;
        POLYGON 3.215 2.93 6.495 2.93 6.495 4.13 8.105 4.13 8.105 1.925 8.335 1.925 8.335 4.36 6.265 4.36 6.265 3.16 3.785 3.16 3.785 4.2 3.555 4.2 3.555 3.16 2.985 3.16 2.985 0.85 3.89 0.85 3.89 1.08 3.215 1.08  ;
        POLYGON 7.645 0.795 7.875 0.795 7.875 1.465 8.795 1.465 8.795 1.98 9.39 1.98 9.39 2.21 8.565 2.21 8.565 1.695 7.875 1.695 7.875 3.9 7.645 3.9  ;
        POLYGON 10.615 2.94 11.455 2.94 11.455 3.9 11.225 3.9 11.225 3.17 10.385 3.17 10.385 0.85 11.33 0.85 11.33 1.08 10.615 1.08  ;
        POLYGON 9.685 0.795 10.115 0.795 10.115 4.13 11.785 4.13 11.785 2.93 12.685 2.93 12.685 1.925 12.915 1.925 12.915 3.16 12.015 3.16 12.015 4.36 9.685 4.36  ;
        POLYGON 13.285 0.795 13.515 0.795 13.515 1.29 14.235 1.29 14.235 1.98 15.74 1.98 15.74 2.21 14.235 2.21 14.235 4.2 14.005 4.2 14.005 1.52 13.285 1.52  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.64 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.35 1.77 11.675 1.77 11.675 2.71 11.35 2.71  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.77 2.65 1.77 2.65 2.71 2.39 2.71  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4716 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.275 0.815 16.65 0.815 16.65 4.21 16.275 4.21  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.435 4.59 1.435 3.4 1.665 3.4 1.665 4.59 2.715 4.59 5.805 4.59 5.805 3.4 6.035 3.4 6.035 4.59 8.345 4.59 8.625 4.59 8.625 3.4 8.855 3.4 8.855 4.59 9.35 4.59 12.025 4.59 12.025 3.4 12.255 3.4 12.255 4.59 12.695 4.59 15.255 4.59 15.255 3.4 15.485 3.4 15.485 4.59 15.98 4.59 17.295 4.59 17.295 3.4 17.525 3.4 17.525 4.59 17.92 4.59 17.92 5.49 15.98 5.49 12.695 5.49 9.35 5.49 8.345 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.675 0.45 17.675 1.625 17.445 1.625 17.445 0.45 15.435 0.45 15.435 1.625 15.205 1.625 15.205 0.45 14.395 0.45 14.395 1.155 14.165 1.155 14.165 0.45 12.155 0.45 12.155 1.155 11.925 1.155 11.925 0.45 8.755 0.45 8.755 1.155 8.525 1.155 8.525 0.45 5.795 0.45 5.795 1.155 5.565 1.155 5.565 0.45 1.65 0.45 1.65 1.1 1.31 1.1 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.815 0.475 0.815 0.475 1.31 1.16 1.31 1.16 1.33 2.065 1.33 2.065 0.815 2.715 0.815 2.715 1.155 2.295 1.155 2.295 1.56 1.065 1.56 1.065 1.54 0.245 1.54  ;
        POLYGON 3.39 1.845 6.685 1.845 6.685 0.815 7.055 0.815 7.055 3.9 6.825 3.9 6.825 2.075 4.775 2.075 4.775 2.71 4.435 2.71 4.435 2.075 3.39 2.075  ;
        POLYGON 3.16 2.835 4.24 2.835 4.24 2.94 6.495 2.94 6.495 4.13 8.115 4.13 8.115 1.885 8.345 1.885 8.345 4.36 6.265 4.36 6.265 3.17 4.275 3.17 4.275 4.21 4.045 4.21 4.045 3.065 2.93 3.065 2.93 1.385 3.605 1.385 3.605 0.815 3.835 0.815 3.835 1.615 3.16 1.615  ;
        POLYGON 7.405 0.815 7.635 0.815 7.635 1.425 8.805 1.425 8.805 1.94 9.35 1.94 9.35 2.17 8.575 2.17 8.575 1.655 7.835 1.655 7.835 3.9 7.405 3.9  ;
        POLYGON 10.535 2.91 11.235 2.91 11.235 3.72 11.005 3.72 11.005 3.14 10.305 3.14 10.305 1.31 11.09 1.31 11.09 1.54 10.535 1.54  ;
        POLYGON 9.645 0.815 9.875 0.815 9.875 3.98 11.565 3.98 11.565 2.94 12.465 2.94 12.465 2.415 12.695 2.415 12.695 3.17 11.795 3.17 11.795 4.21 9.645 4.21  ;
        POLYGON 12.99 1.31 13.33 1.31 13.33 1.33 14.015 1.33 14.015 1.94 15.98 1.94 15.98 2.17 14.015 2.17 14.015 4.21 13.785 4.21 13.785 1.56 12.99 1.56  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.16 BY 5.04 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.64 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.35 1.77 11.61 1.77 11.61 2.71 11.35 2.71  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.345 1.82 2.65 1.82 2.65 3.27 2.345 3.27  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.03 2.69 17.51 2.69 18.07 2.69 18.07 1.6 16.03 1.6 16.03 0.79 16.31 0.79 16.31 1.3 18.32 1.3 18.32 0.79 18.55 0.79 18.55 3.96 18.07 3.96 18.07 2.92 17.51 2.92 16.26 2.92 16.26 3.96 16.03 3.96  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.325 4.59 1.325 3.15 1.555 3.15 1.555 4.59 2.715 4.59 5.82 4.59 5.82 3.15 6.05 3.15 6.05 4.59 8.25 4.59 8.58 4.59 8.58 3.15 8.81 3.15 8.81 4.59 9.305 4.59 12.08 4.59 12.08 3.785 12.31 3.785 12.31 4.59 12.75 4.59 15.01 4.59 15.01 3.15 15.24 3.15 15.24 4.59 17.05 4.59 17.05 3.15 17.28 3.15 17.28 4.59 17.51 4.59 19.09 4.59 19.09 3.15 19.32 3.15 19.32 4.59 20.16 4.59 20.16 5.49 17.51 5.49 12.75 5.49 9.305 5.49 8.25 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.16 -0.45 20.16 0.45 19.67 0.45 19.67 1.6 19.44 1.6 19.44 0.45 17.43 0.45 17.43 1.07 17.2 1.07 17.2 0.45 15.19 0.45 15.19 1.6 14.96 1.6 14.96 0.45 14.45 0.45 14.45 1.13 14.22 1.13 14.22 0.45 12.21 0.45 12.21 1.13 11.98 1.13 11.98 0.45 8.81 0.45 8.81 1.13 8.58 1.13 8.58 0.45 5.81 0.45 5.81 1.13 5.58 1.13 5.58 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 1.305 2.485 1.305 2.485 0.79 2.715 0.79 2.715 1.535 0.245 1.535  ;
        POLYGON 3.405 1.845 6.7 1.845 6.7 0.79 7.07 0.79 7.07 3.9 6.84 3.9 6.84 2.075 4.81 2.075 4.81 2.46 4.47 2.46 4.47 2.075 3.405 2.075  ;
        POLYGON 3.175 2.565 4.265 2.565 4.265 2.69 6.51 2.69 6.51 4.13 8.02 4.13 8.02 1.82 8.25 1.82 8.25 4.36 6.28 4.36 6.28 2.92 4.29 2.92 4.29 3.96 4.06 3.96 4.06 2.795 2.945 2.795 2.945 1.385 3.62 1.385 3.62 0.79 3.85 0.79 3.85 1.615 3.175 1.615  ;
        POLYGON 7.46 0.79 7.69 0.79 7.69 1.36 8.71 1.36 8.71 1.875 9.305 1.875 9.305 2.105 8.48 2.105 8.48 1.59 7.79 1.59 7.79 3.9 7.46 3.9  ;
        POLYGON 10.36 1.23 11.09 1.23 11.09 2.935 11.29 2.935 11.29 3.275 10.86 3.275 10.86 1.46 10.59 1.46 10.59 2.2 10.36 2.2  ;
        POLYGON 9.6 0.79 9.93 0.79 9.93 3.505 11.63 3.505 11.63 3.325 12.52 3.325 12.52 2.475 12.75 2.475 12.75 3.555 11.855 3.555 11.855 3.735 9.83 3.735 9.83 3.96 9.6 3.96  ;
        POLYGON 13.045 1.285 13.385 1.285 13.385 1.305 14.07 1.305 14.07 1.98 17.51 1.98 17.51 2.32 14.07 2.32 14.07 3.96 13.84 3.96 13.84 1.535 13.045 1.535  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.12 BY 5.04 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.22 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.23 1.77 10.49 1.77 10.49 2.71 10.23 2.71  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.255 1.77 2.255 2.71 1.83 2.71  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.21 0.41 1.21 0.41 2.27 1.19 2.27 1.19 2.5 0.15 2.5  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2452 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.15 0.695 14.61 0.695 14.61 3.685 14.15 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.21 4.59 13.915 4.59 15.12 4.59 15.12 5.49 13.915 5.49 2.935 5.49 0 5.49 0 4.59 0.845 4.59 0.845 3.435 1.075 3.435 1.075 4.59 2.935 4.59 6.025 4.59 6.025 3.91 6.255 3.91 6.255 4.59 8.98 4.59 8.98 3.895 11.2 3.895 11.2 4.005 13.01 4.005 13.01 3.425 13.24 3.425 13.24 4.235 9.21 4.235  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.12 -0.45 15.12 0.45 13.49 0.45 13.49 1.015 13.26 1.015 13.26 0.45 9.49 0.45 9.49 1.035 9.26 1.035 9.26 0.45 6.015 0.45 6.015 1.13 5.785 1.13 5.785 0.45 1.87 0.45 1.87 1.075 1.53 1.075 1.53 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.75 0.87 0.75 0.87 1.305 2.705 1.305 2.705 0.79 2.935 0.79 2.935 1.535 0.64 1.535 0.64 0.98 0.19 0.98  ;
        POLYGON 3.665 1.79 3.895 1.79 3.895 2.485 4.99 2.485 4.99 2.715 3.665 2.715  ;
        POLYGON 3.435 2.945 5.22 2.945 5.22 1.755 6.37 1.755 6.37 2.27 6.75 2.27 6.75 2.5 6.14 2.5 6.14 1.985 5.45 1.985 5.45 3.175 3.595 3.175 3.595 4.245 3.205 4.245 3.205 0.845 4.11 0.845 4.11 1.075 3.435 1.075  ;
        POLYGON 7.565 2.375 8.14 2.375 8.14 0.695 8.475 0.695 8.475 3.18 8.135 3.18 8.135 2.605 7.565 2.605  ;
        POLYGON 8.715 2.27 9.77 2.27 9.77 0.75 10.665 0.75 10.665 0.98 10 0.98 10 2.95 10.515 2.95 10.515 3.18 9.77 3.18 9.77 2.5 8.715 2.5  ;
        POLYGON 5.68 2.215 5.91 2.215 5.91 3.41 6.98 3.41 6.98 1.13 6.905 1.13 6.905 0.79 7.21 0.79 7.21 3.41 10.745 3.41 10.745 2.27 12.555 2.27 12.555 2.5 10.975 2.5 10.975 3.64 7.275 3.64 7.275 4.245 7.045 4.245 7.045 3.64 5.68 3.64  ;
        POLYGON 11.99 2.875 12.785 2.875 12.785 1.035 11.1 1.035 11.1 0.695 13.015 0.695 13.015 2.27 13.915 2.27 13.915 2.5 13.015 2.5 13.015 3.105 12.22 3.105 12.22 3.685 11.99 3.685  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.625 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.23 1.21 10.425 1.21 10.49 1.21 10.49 2.405 10.425 2.405 10.23 2.405  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 1.77 2.09 1.77 2.09 2.35 1.21 2.35  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4716 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.59 2.89 13.94 2.89 13.94 1.59 13.59 1.59 13.59 1.21 13.94 1.21 13.94 0.79 14.2 0.79 14.2 3.685 13.59 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.95 4.59 13.49 4.59 15.68 4.59 15.68 5.49 13.49 5.49 2.715 5.49 0 5.49 0 4.59 0.695 4.59 0.695 3.44 0.925 3.44 0.925 4.59 2.715 4.59 5.805 4.59 5.805 3.85 6.035 3.85 6.035 4.59 8.72 4.59 8.72 3.85 11.14 3.85 11.14 4.02 12.95 4.02 12.95 3.44 13.18 3.44 13.18 4.02 13.49 4.02 14.99 4.02 14.99 3.44 15.22 3.44 15.22 4.25 13.49 4.25 8.95 4.25  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 15.29 0.45 15.29 1.43 15.06 1.43 15.06 0.45 13.05 0.45 13.05 1.43 12.82 1.43 12.82 0.45 9.25 0.45 9.25 1.13 9.02 1.13 9.02 0.45 5.85 0.45 5.85 1.13 5.62 1.13 5.62 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 1.305 2.485 1.305 2.485 0.79 2.715 0.79 2.715 1.535 0.245 1.535  ;
        POLYGON 3.445 1.79 3.675 1.79 3.675 2.485 4.77 2.485 4.77 2.715 3.445 2.715  ;
        POLYGON 3.215 2.945 5 2.945 5 1.605 6.345 1.605 6.345 2.35 6.005 2.35 6.005 1.835 5.23 1.835 5.23 3.175 3.785 3.175 3.785 4.25 3.555 4.25 3.555 3.175 2.985 3.175 2.985 0.845 3.89 0.845 3.89 1.075 3.215 1.075  ;
        POLYGON 7.4 0.845 8.185 0.845 8.185 1.075 7.63 1.075 7.63 2.93 7.985 2.93 7.985 3.16 7.4 3.16  ;
        POLYGON 8.225 2.12 9.685 2.12 9.685 0.75 10.425 0.75 10.425 0.98 9.915 0.98 9.915 2.93 10.025 2.93 10.025 3.16 9.685 3.16 9.685 2.35 8.225 2.35  ;
        POLYGON 5.46 2.065 5.69 2.065 5.69 3.39 6.74 3.39 6.74 0.79 6.97 0.79 6.97 3.39 11.47 3.39 11.47 2.12 12.425 2.12 12.425 2.35 11.7 2.35 11.7 3.62 7.055 3.62 7.055 4.25 6.825 4.25 6.825 3.62 5.46 3.62  ;
        POLYGON 11.93 2.875 12.655 2.875 12.655 1.89 10.86 1.89 10.86 0.79 11.09 0.79 11.09 1.66 12.885 1.66 12.885 2.065 13.49 2.065 13.49 2.405 12.885 2.405 12.885 3.105 12.16 3.105 12.16 3.685 11.93 3.685  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.625 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.23 1.77 10.315 1.77 10.49 1.77 10.49 2.71 10.315 2.71 10.23 2.71  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.175 2.09 2.175 2.09 2.405 0.97 2.405 0.97 2.71 0.71 2.71  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.415 1.77 0.415 2.71 0.15 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.885 2.875 15.37 2.875 15.955 2.875 15.955 1.745 13.885 1.745 13.885 0.795 14.115 0.795 14.115 1.515 15.77 1.515 15.77 0.71 16.355 0.71 16.355 3.685 15.955 3.685 15.955 3.105 15.37 3.105 14.145 3.105 14.145 3.685 13.885 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.125 4.59 15.37 4.59 17.92 4.59 17.92 5.49 15.37 5.49 2.715 5.49 0 5.49 0 4.59 0.625 4.59 0.625 3.44 0.855 3.44 0.855 4.59 2.715 4.59 5.805 4.59 5.805 3.855 6.035 3.855 6.035 4.59 8.865 4.59 8.865 3.855 9.095 3.855 9.095 4.59 10.855 4.59 10.855 3.855 11.085 3.855 11.085 4.59 12.895 4.59 12.895 3.44 13.125 3.44 13.125 4.02 14.935 4.02 14.935 3.44 15.165 3.44 15.165 4.02 15.37 4.02 16.975 4.02 16.975 3.44 17.205 3.44 17.205 4.25 15.37 4.25 13.125 4.25  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.475 0.45 17.475 1.485 17.245 1.485 17.245 0.45 15.235 0.45 15.235 1.035 15.005 1.035 15.005 0.45 12.995 0.45 12.995 1.485 12.765 1.485 12.765 0.45 9.195 0.45 9.195 1.135 8.965 1.135 8.965 0.45 5.795 0.45 5.795 1.135 5.565 1.135 5.565 0.45 1.65 0.45 1.65 1.08 1.31 1.08 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.795 0.475 0.795 0.475 1.31 2.485 1.31 2.485 0.795 2.715 0.795 2.715 1.54 0.245 1.54  ;
        POLYGON 3.445 1.79 4.715 1.79 4.715 2.77 4.485 2.77 4.485 2.13 3.445 2.13  ;
        POLYGON 3.215 2.82 4.26 2.82 4.26 3 4.945 3 4.945 1.66 6.095 1.66 6.095 2.175 6.53 2.175 6.53 2.405 5.865 2.405 5.865 1.89 5.175 1.89 5.175 3.23 4.265 3.23 4.265 4.25 4.035 4.25 4.035 3.05 2.985 3.05 2.985 0.85 3.89 0.85 3.89 1.08 3.215 1.08  ;
        POLYGON 7.345 2.12 7.845 2.12 7.845 0.795 8.13 0.795 8.13 3.16 7.79 3.16 7.79 2.46 7.345 2.46  ;
        POLYGON 8.37 2.175 9.77 2.175 9.77 1.31 10.085 1.31 10.085 0.795 10.315 0.795 10.315 1.54 10 1.54 10 2.935 10.17 2.935 10.17 3.165 9.77 3.165 9.77 2.405 8.37 2.405  ;
        POLYGON 5.405 2.12 5.635 2.12 5.635 3.395 6.76 3.395 6.76 1.135 6.685 1.135 6.685 0.795 6.99 0.795 6.99 3.395 11.415 3.395 11.415 2.175 12.6 2.175 12.6 2.405 11.645 2.405 11.645 3.625 7.055 3.625 7.055 4.25 6.825 4.25 6.825 3.625 5.405 3.625  ;
        POLYGON 11.875 2.875 12.83 2.875 12.83 1.945 10.805 1.945 10.805 0.795 11.035 0.795 11.035 1.715 13.06 1.715 13.06 1.975 15.37 1.975 15.37 2.315 13.06 2.315 13.06 3.105 12.105 3.105 12.105 3.685 11.875 3.685  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.24 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.21 1.015 1.21 1.015 2.3 1.07 2.3 1.07 2.53 0.71 2.53  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 0.68 1.595 0.68 1.595 4.36 1.365 4.36 1.365 2.15 1.27 2.15  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 2.24 4.59 2.24 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.24 -0.45 2.24 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 3.36 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 1.91 2.27 1.91 2.71 0.63 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9155 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.395 3.45 2.14 3.45 2.14 1.85 1.83 1.85 1.83 1.49 1.395 1.49 1.395 0.68 1.625 0.68 1.625 1.21 2.285 1.21 2.285 1.67 2.37 1.67 2.37 3.83 1.625 3.83 1.625 4.36 1.395 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.6 4.59 2.6 3.55 2.83 3.55 2.83 4.59 3.36 4.59 3.36 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 3.36 -0.45 3.36 0.45 2.745 0.45 2.745 1.49 2.515 1.49 2.515 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.121 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 2.27 2.16 2.27 2.16 2.71 0.41 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.207 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 2.39 3.09 2.39 1.95 1.365 1.95 1.365 0.68 1.595 0.68 1.595 1.72 3.605 1.72 3.605 0.68 3.835 0.68 3.835 1.95 2.805 1.95 2.805 3.09 3.735 3.09 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.48 4.59 4.48 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_3
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.58 2.27 2.33 2.27 2.33 2.65 0.58 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.12 3.335 3.12 3.335 1.89 1.365 1.89 1.365 0.68 1.595 0.68 1.595 1.66 3.605 1.66 3.605 0.68 3.835 0.68 3.835 4.36 3.505 4.36 3.505 3.35 1.595 3.35 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.58 2.615 3.58 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 5.6 4.59 5.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.955 0.45 4.955 1.43 4.725 1.43 4.725 0.45 2.715 0.45 2.715 1.43 2.485 1.43 2.485 0.45 0.475 0.45 0.475 1.43 0.245 1.43 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.656 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.265 4.26 2.265 4.26 2.645 0.63 2.645  ;
        POLYGON 5.36 2.215 8.88 2.215 8.88 2.65 5.36 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 4.63 3.09 4.63 1.985 1.365 1.985 1.365 0.68 1.595 0.68 1.595 1.755 3.575 1.755 3.575 0.68 3.835 0.68 3.835 1.755 5.845 1.755 5.845 0.68 6.075 0.68 6.075 1.755 8.085 1.755 8.085 0.68 8.315 0.68 8.315 1.985 5.13 1.985 5.13 3.09 8.215 3.09 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 10.08 4.59 10.08 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.165 4.725 1.165 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_8
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 20.484 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.18 2.27 5.69 2.27 5.69 2.65 0.18 2.65  ;
        POLYGON 7.6 2.215 13 2.215 13 2.65 7.6 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.926 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 6.755 3.09 6.755 1.95 1.365 1.95 1.365 0.68 1.625 0.68 1.625 1.72 3.605 1.72 3.605 0.68 3.835 0.68 3.835 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 1.72 8.085 1.72 8.085 0.68 8.315 0.68 8.315 1.72 10.325 1.72 10.325 0.68 10.555 0.68 10.555 1.72 12.565 1.72 12.565 0.68 12.795 0.68 12.795 1.95 7.37 1.95 7.37 3.09 12.695 3.09 12.695 4.36 12.465 4.36 12.465 3.32 10.455 3.32 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 14.56 4.59 14.56 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_12
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 27.312 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.215 7.965 2.215 7.965 2.65 0.685 2.65  ;
        POLYGON 9.225 2.215 16.505 2.215 16.505 2.65 9.225 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.568 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.98 8.195 2.98 8.195 1.95 1.365 1.95 1.365 0.68 1.625 0.68 1.625 1.72 3.605 1.72 3.605 0.68 3.835 0.68 3.835 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 1.72 8.085 1.72 8.085 0.68 8.315 0.68 8.315 1.72 10.325 1.72 10.325 0.68 10.555 0.68 10.555 1.72 12.565 1.72 12.565 0.68 12.795 0.68 12.795 1.72 14.805 1.72 14.805 0.68 15.035 0.68 15.035 1.72 17.045 1.72 17.045 0.68 17.275 0.68 17.275 1.95 8.995 1.95 8.995 2.95 17.175 2.95 17.175 4.36 16.945 4.36 16.945 3.18 14.935 3.18 14.935 4.36 14.705 4.36 14.705 3.18 12.695 3.18 12.695 4.36 12.465 4.36 12.465 3.18 10.455 3.18 10.455 4.36 10.225 4.36 10.225 3.18 8.31 3.18 8.31 4.36 8.08 4.36 8.08 3.21 5.975 3.21 5.975 4.36 5.745 4.36 5.745 3.21 3.735 3.21 3.735 4.36 3.505 4.36 3.505 3.21 1.595 3.21 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 19.04 4.59 19.04 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 18.395 0.45 18.395 1.49 18.165 1.49 18.165 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_16
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 34.14 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 9.9 2.27 9.9 2.65 0.63 2.65  ;
        POLYGON 11.11 2.27 20.38 2.27 20.38 2.65 11.11 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 18.21 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 10.13 3.09 10.13 1.95 1.335 1.95 1.335 0.68 1.595 0.68 1.595 1.72 3.605 1.72 3.605 0.68 3.835 0.68 3.835 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 1.72 8.085 1.72 8.085 0.68 8.315 0.68 8.315 1.72 10.325 1.72 10.325 0.68 10.555 0.68 10.555 1.72 12.565 1.72 12.565 0.68 12.795 0.68 12.795 1.72 14.805 1.72 14.805 0.68 15.035 0.68 15.035 1.72 17.045 1.72 17.045 0.68 17.275 0.68 17.275 1.72 19.285 1.72 19.285 0.68 19.515 0.68 19.515 1.72 21.525 1.72 21.525 0.68 21.755 0.68 21.755 1.95 10.88 1.95 10.88 3.09 21.655 3.09 21.655 4.36 21.425 4.36 21.425 3.32 19.415 3.32 19.415 4.36 19.185 4.36 19.185 3.32 17.175 3.32 17.175 4.36 16.945 4.36 16.945 3.32 14.935 3.32 14.935 4.36 14.705 4.36 14.705 3.32 12.695 3.32 12.695 4.36 12.465 4.36 12.465 3.32 10.455 3.32 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 20.305 4.59 20.305 3.55 20.535 3.55 20.535 4.59 22.545 4.59 22.545 3.55 22.775 3.55 22.775 4.59 23.52 4.59 23.52 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 22.875 0.45 22.875 1.49 22.645 1.49 22.645 0.45 20.635 0.45 20.635 1.49 20.405 1.49 20.405 0.45 18.395 0.45 18.395 1.49 18.165 1.49 18.165 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_20
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.698 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.015 0.97 2.015 0.97 2.71 0.15 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.849 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.505 1.77 8.81 1.77 8.81 2.71 8.505 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.3728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 1.14 4.84 1.14 4.84 1.77 4.89 1.77 4.89 3.9 4.61 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.48 1.495 3.48 1.495 4.59 5.68 4.59 5.68 3.86 5.91 3.86 5.91 4.59 6.795 4.59 7.585 4.59 7.585 3.48 7.815 3.48 7.815 4.59 9.33 4.59 9.52 4.59 9.52 5.49 9.33 5.49 6.795 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 7.815 0.45 7.815 1.48 7.585 1.48 7.585 0.45 5.96 0.45 5.96 1.165 5.73 1.165 5.73 0.45 1.84 0.45 1.84 1.48 1.61 1.48 1.61 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.02 2.105 3.02 2.105 2.245 1.2 2.245 1.2 1.82 1.095 1.82 1.095 1.425 0.19 1.425 0.19 1.195 1.325 1.195 1.325 1.625 1.43 1.625 1.43 2.015 2.335 2.015 2.335 3.02 3.06 3.02 3.06 3.25 0.475 3.25 0.475 4.29 0.245 4.29  ;
        POLYGON 2.675 1.195 3.355 1.195 3.355 0.68 5.3 0.68 5.3 1.395 6.465 1.395 6.465 1.14 6.695 1.14 6.695 1.625 5.375 1.625 5.375 2.17 5.145 2.17 5.145 1.565 5.07 1.565 5.07 0.91 3.585 0.91 3.585 3.82 3.355 3.82 3.355 1.425 2.675 1.425  ;
        POLYGON 2.335 3.48 2.565 3.48 2.565 4.13 3.85 4.13 3.85 1.14 4.08 1.14 4.08 4.13 5.12 4.13 5.12 2.43 5.415 2.43 5.415 3.4 6.795 3.4 6.795 4.29 6.565 4.29 6.565 3.63 5.35 3.63 5.35 4.36 2.335 4.36  ;
        POLYGON 7.09 2.015 8.045 2.015 8.045 1.195 9.33 1.195 9.33 1.425 8.275 1.425 8.275 3.15 9.175 3.15 9.175 4.29 8.945 4.29 8.945 3.38 8.045 3.38 8.045 2.245 7.09 2.245  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.99 1.77 8.46 1.77 8.46 2.71 7.99 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.62 0.68 6.85 0.68 6.85 1.21 7.13 1.21 7.13 2.71 7 2.71 7 3.75 6.77 3.75 6.77 1.49 6.62 1.49  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.37 4.59 1.37 3.4 1.6 3.4 1.6 4.59 5.75 4.59 5.75 4.35 5.98 4.35 5.98 4.59 7.79 4.59 7.79 3.4 8.02 3.4 8.02 4.59 9.09 4.59 9.52 4.59 9.52 5.49 9.09 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 7.97 0.45 7.97 1.49 7.74 1.49 7.74 0.45 5.73 0.45 5.73 1.02 5.5 1.02 5.5 0.45 1.65 0.45 1.65 1.02 1.42 1.02 1.42 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.35 2.94 1.86 2.94 1.86 1.49 0.3 1.49 0.3 0.68 0.53 0.68 0.53 1.26 2.09 1.26 2.09 2.47 3.625 2.47 3.625 3.17 0.58 3.17 0.58 4.21 0.35 4.21  ;
        POLYGON 2.54 0.68 5.265 0.68 5.265 1.25 6.39 1.25 6.39 2.11 6.16 2.11 6.16 1.48 5.035 1.48 5.035 1.085 3.43 1.085 3.43 2.01 4.15 2.01 4.15 3.9 3.92 3.9 3.92 2.24 3.2 2.24 3.2 1.49 2.54 1.49  ;
        POLYGON 2.9 3.4 3.13 3.4 3.13 4.13 4.585 4.13 4.585 1.78 3.66 1.78 3.66 1.315 3.89 1.315 3.89 1.55 4.815 1.55 4.815 1.99 5.93 1.99 5.93 2.465 6.475 2.465 6.475 2.695 5.7 2.695 5.7 2.22 4.96 2.22 4.96 4.36 2.9 4.36  ;
        POLYGON 5.24 2.45 5.47 2.45 5.47 2.925 6.395 2.925 6.395 3.98 7.33 3.98 7.33 2.94 8.86 2.94 8.86 0.68 9.09 0.68 9.09 4.21 8.81 4.21 8.81 3.17 7.56 3.17 7.56 4.21 6.165 4.21 6.165 3.155 5.24 3.155  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.88 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 1.77 5.645 1.77 5.645 2.71 5.19 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9952 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.465 2.965 11.365 2.965 12.03 2.965 12.265 2.965 12.265 1.6 10.025 1.6 10.025 0.79 10.255 0.79 10.255 1.37 12.265 1.37 12.265 0.84 12.495 0.84 12.495 3.195 12.03 3.195 11.735 3.195 11.735 4.21 11.505 4.21 11.505 3.195 11.365 3.195 9.93 3.195 9.93 4.21 9.465 4.21  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.37 4.59 1.37 3.845 1.6 3.845 1.6 4.59 6.045 4.59 6.045 4.28 6.275 4.28 6.275 4.59 8.265 4.59 8.265 3.4 8.495 3.4 8.495 4.59 10.485 4.59 10.485 3.88 10.715 3.88 10.715 4.59 11.365 4.59 12.03 4.59 12.88 4.59 12.88 5.49 12.03 5.49 11.365 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.88 -0.45 12.88 0.45 11.375 0.45 11.375 1.02 11.145 1.02 11.145 0.45 8.955 0.45 8.955 1.16 8.725 1.16 8.725 0.45 6.575 0.45 6.575 0.62 6.235 0.62 6.235 0.45 1.65 0.45 1.65 1.02 1.42 1.02 1.42 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.35 2.94 3.335 2.94 3.335 2.06 1.2 2.06 1.2 1.54 0.3 1.54 0.3 0.68 0.53 0.68 0.53 1.31 1.43 1.31 1.43 1.83 3.565 1.83 3.565 3.17 0.58 3.17 0.58 4.21 0.35 4.21  ;
        POLYGON 5.025 2.94 6.75 2.94 6.75 1.54 4.92 1.54 4.92 1.31 7.09 1.31 7.09 2.06 6.98 2.06 6.98 3.17 5.255 3.17 5.255 3.75 5.025 3.75  ;
        POLYGON 2.895 3.4 3.125 3.4 3.125 3.98 4.375 3.98 4.375 1.655 4.255 1.655 4.255 1.315 4.605 1.315 4.605 3.98 5.605 3.98 5.605 3.82 7.245 3.82 7.245 2.505 11.365 2.505 11.365 2.735 7.475 2.735 7.475 4.05 5.825 4.05 5.825 4.21 2.895 4.21  ;
        POLYGON 2.54 0.68 2.77 0.68 2.77 0.85 7.835 0.85 7.835 1.83 12.03 1.83 12.03 2.06 7.605 2.06 7.605 1.08 4.025 1.08 4.025 2.94 4.145 2.94 4.145 3.75 3.795 3.75 3.795 1.49 2.54 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_3
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 13.44 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 1.02 1.77 1.02 2.06 0.41 2.06 0.41 2.71 0.15 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.83 6.07 1.83 6.07 2.65 5.13 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.2448 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.11 2.965 11.075 2.965 11.585 2.965 11.585 1.62 9.18 1.62 9.18 0.73 9.63 0.73 9.63 1.39 11.64 1.39 11.64 0.73 11.87 0.73 11.87 3.9 11.19 3.9 11.19 3.31 11.075 3.31 9.41 3.31 9.41 3.9 9.11 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.845 1.545 3.845 1.545 4.59 6.04 4.59 6.04 3.8 6.27 3.8 6.27 4.59 8.13 4.59 8.13 3.88 8.36 3.88 8.36 4.59 10.17 4.59 10.17 3.88 10.4 3.88 10.4 4.59 11.075 4.59 12.21 4.59 12.21 3.09 12.44 3.09 12.44 4.59 13.44 4.59 13.44 5.49 11.075 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 13.44 -0.45 13.44 0.45 12.99 0.45 12.99 1.54 12.76 1.54 12.76 0.45 10.75 0.45 10.75 1.16 10.52 1.16 10.52 0.45 8.51 0.45 8.51 0.69 8.28 0.69 8.28 0.45 6.325 0.45 6.325 0.635 5.985 0.635 5.985 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 3.09 1.25 3.09 1.25 1.54 0.245 1.54 0.245 0.73 0.475 0.73 0.475 1.31 1.48 1.31 1.48 1.83 2.09 1.83 2.09 2.29 3.595 2.29 3.595 2.755 3.365 2.755 3.365 2.52 1.86 2.52 1.86 2.06 1.48 2.06 1.48 3.32 0.525 3.32 0.525 3.9 0.295 3.9  ;
        POLYGON 5.02 2.88 6.53 2.88 6.53 1.595 4.865 1.595 4.865 1.365 6.76 1.365 6.76 3.11 5.25 3.11 5.25 3.9 5.02 3.9  ;
        POLYGON 2.485 0.73 3.315 0.73 3.315 0.905 7.445 0.905 7.445 1.04 8.95 1.04 8.95 1.85 10.265 1.85 10.265 2.11 8.72 2.11 8.72 1.27 7.235 1.27 7.235 1.135 3.32 1.135 3.32 1.83 4.175 1.83 4.175 3.9 3.945 3.9 3.945 2.06 3.09 2.06 3.09 0.96 2.715 0.96 2.715 1.54 2.485 1.54  ;
        POLYGON 2.925 3.09 3.155 3.09 3.155 4.13 4.405 4.13 4.405 1.6 3.55 1.6 3.55 1.37 4.635 1.37 4.635 4.13 5.58 4.13 5.58 3.34 7.115 3.34 7.115 2.505 11.075 2.505 11.075 2.735 7.345 2.735 7.345 4.15 7.11 4.15 7.11 3.57 5.81 3.57 5.81 4.36 2.925 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.72 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.77 1.555 1.77 1.555 2.71 1.27 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 2.33 5.45 2.33 5.45 3.27 5.165 3.27  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.6696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.215 2.925 17.195 2.925 17.535 2.925 18.315 2.925 18.315 1.595 12.165 1.595 12.165 0.68 12.395 0.68 12.395 1.21 14.405 1.21 14.405 0.68 14.635 0.68 14.635 1.215 16.645 1.215 16.645 0.68 16.875 0.68 16.875 1.21 18.885 1.21 18.885 0.68 19.115 0.68 19.115 1.595 18.805 1.595 18.805 4.195 18.335 4.195 18.335 3.155 17.535 3.155 17.195 3.155 16.525 3.155 16.525 4.195 16.295 4.195 16.295 3.155 14.485 3.155 14.485 4.19 14.255 4.19 14.255 3.155 12.455 3.155 12.455 4.19 12.215 4.19  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.905 4.59 1.905 3.42 2.135 3.42 2.135 4.59 4.675 4.59 4.675 4.35 4.905 4.35 4.905 4.59 6.715 4.59 6.715 4.35 6.945 4.35 6.945 4.59 8.755 4.59 8.755 3.38 8.985 3.38 8.985 4.59 10.995 4.59 10.995 3.88 11.225 3.88 11.225 4.59 13.235 4.59 13.235 3.385 13.465 3.385 13.465 4.59 15.275 4.59 15.275 3.385 15.505 3.385 15.505 4.59 17.195 4.59 17.315 4.59 17.315 3.385 17.535 3.385 17.545 3.385 17.545 4.59 19.355 4.59 19.355 3.38 19.585 3.38 19.585 4.59 20.72 4.59 20.72 5.49 17.535 5.49 17.195 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.72 -0.45 20.72 0.45 20.235 0.45 20.235 1.49 20.005 1.49 20.005 0.45 17.995 0.45 17.995 0.98 17.765 0.98 17.765 0.45 15.755 0.45 15.755 0.98 15.525 0.98 15.525 0.45 13.515 0.45 13.515 0.98 13.285 0.98 13.285 0.45 11.275 0.45 11.275 1.49 11.045 1.49 11.045 0.45 9.035 0.45 9.035 1.49 8.805 1.49 8.805 0.45 6.85 0.45 6.85 0.635 6.51 0.635 6.51 0.45 4.61 0.45 4.61 0.635 4.27 0.635 4.27 0.45 1.595 0.45 1.595 1.02 1.365 1.02 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.885 2.94 2.63 2.94 2.63 2.11 1.805 2.11 1.805 1.49 0.245 1.49 0.245 0.68 0.475 0.68 0.475 1.26 2.035 1.26 2.035 1.88 2.86 1.88 2.86 2.425 3.65 2.425 3.65 3.15 2.725 3.15 2.725 3.17 1.115 3.17 1.115 4.19 0.885 4.19  ;
        POLYGON 5.695 2.48 7.155 2.48 7.155 1.595 5.39 1.595 5.39 1.365 7.385 1.365 7.385 2.71 5.925 2.71 5.925 3.66 5.695 3.66  ;
        POLYGON 2.925 3.38 3.155 3.38 3.155 3.89 4.405 3.89 4.405 1.595 3.55 1.595 3.55 1.365 4.635 1.365 4.635 3.89 7.735 3.89 7.735 2.405 17.195 2.405 17.195 2.695 10.105 2.695 10.105 4.19 9.875 4.19 9.875 2.695 7.965 2.695 7.965 4.19 7.735 4.19 7.735 4.12 2.925 4.12  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.905 7.63 0.905 7.63 0.855 7.975 0.855 7.975 1.825 9.925 1.825 9.925 0.84 10.155 0.84 10.155 1.825 17.535 1.825 17.535 2.055 7.745 2.055 7.745 1.135 3.32 1.135 3.32 1.825 4.175 1.825 4.175 3.66 3.945 3.66 3.945 2.055 3.09 2.055 3.09 1.49 2.485 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_8
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 29.12 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.076 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.57 1.785 6.01 1.785 6.01 3.27 5.57 3.27  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.2744 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.14 3.01 25.57 3.01 25.94 3.01 26.45 3.01 26.45 1.595 16.09 1.595 16.09 0.895 27.52 0.895 27.52 1.595 26.98 1.595 26.98 3.01 26.97 3.01 26.97 4.28 26.735 4.28 26.735 3.49 25.94 3.49 25.57 3.49 24.93 3.49 24.93 4.28 24.7 4.28 24.7 3.49 22.89 3.49 22.89 4.28 22.66 4.28 22.66 3.49 20.75 3.49 20.75 4.28 20.52 4.28 20.52 3.49 18.51 3.49 18.51 4.28 18.28 4.28 18.28 3.49 16.37 3.49 16.37 4.28 16.14 4.28  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.83 4.59 1.83 3.47 2.06 3.47 2.06 4.59 6.03 4.59 6.03 4.51 6.26 4.51 6.26 4.59 8.51 4.59 8.51 4.51 8.74 4.51 8.74 4.59 10.77 4.59 10.77 3.95 11 3.95 11 4.59 12.81 4.59 12.81 3.47 13.04 3.47 13.04 4.59 14.92 4.59 14.92 3.88 15.15 3.88 15.15 4.59 17.16 4.59 17.16 3.96 17.39 3.96 17.39 4.59 19.4 4.59 19.4 3.94 19.63 3.94 19.63 4.59 21.64 4.59 21.64 3.94 21.87 3.94 21.87 4.59 23.68 4.59 23.68 3.94 23.91 3.94 23.91 4.59 25.57 4.59 25.72 4.59 25.72 3.94 25.94 3.94 25.95 3.94 25.95 4.59 27.76 4.59 27.76 3.47 27.99 3.47 27.99 4.59 29.12 4.59 29.12 5.49 25.94 5.49 25.57 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 29.12 -0.45 29.12 0.45 28.64 0.45 28.64 1.54 28.41 1.54 28.41 0.45 26.455 0.45 26.455 0.635 26.115 0.635 26.115 0.45 24.215 0.45 24.215 0.635 23.875 0.635 23.875 0.45 21.975 0.45 21.975 0.635 21.635 0.635 21.635 0.45 19.735 0.45 19.735 0.635 19.395 0.635 19.395 0.45 17.495 0.45 17.495 0.635 17.155 0.635 17.155 0.45 15.2 0.45 15.2 1.54 14.97 1.54 14.97 0.45 12.96 0.45 12.96 1.54 12.73 1.54 12.73 0.45 10.72 0.45 10.72 1.54 10.49 1.54 10.49 0.45 8.535 0.45 8.535 0.635 8.195 0.635 8.195 0.45 6.295 0.45 6.295 0.635 5.955 0.635 5.955 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.81 2.94 1.805 2.94 1.805 1.54 0.245 1.54 0.245 0.73 0.475 0.73 0.475 1.31 2.035 1.31 2.035 2.48 3.575 2.48 3.575 3.17 1.04 3.17 1.04 4.28 0.81 4.28  ;
        POLYGON 4.79 3.01 5.02 3.01 5.02 3.59 7.27 3.59 7.27 2.23 8.69 2.23 8.69 1.555 4.835 1.555 4.835 1.325 8.975 1.325 8.975 2.525 7.5 2.525 7.5 3.82 4.79 3.82  ;
        POLYGON 2.85 3.47 3.08 3.47 3.08 4.05 4.33 4.05 4.33 1.595 3.55 1.595 3.55 1.365 4.56 1.365 4.56 4.05 9.75 4.05 9.75 2.505 25.57 2.505 25.57 2.735 14.06 2.735 14.06 4.28 13.83 4.28 13.83 2.735 12.02 2.735 12.02 4.28 11.79 4.28 11.79 2.735 9.98 2.735 9.98 4.28 2.85 4.28  ;
        POLYGON 2.485 0.73 2.715 0.73 2.715 0.865 9.315 0.865 9.315 0.815 9.66 0.815 9.66 1.825 11.61 1.825 11.61 0.84 11.84 0.84 11.84 1.825 13.85 1.825 13.85 0.84 14.08 0.84 14.08 1.825 25.94 1.825 25.94 2.055 9.43 2.055 9.43 1.095 3.32 1.095 3.32 1.825 4.1 1.825 4.1 3.82 3.87 3.82 3.87 2.055 3.09 2.055 3.09 1.095 2.715 1.095 2.715 1.54 2.485 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_12
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 36.96 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.815 1.85 1.155 1.85 1.155 2.275 0.815 2.275  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.768 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.065 2.03 7.71 2.03 7.71 2.605 5.065 2.605  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.3292 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.405 2.965 33.7 2.965 33.73 2.965 34.835 2.965 34.835 1.595 19.405 1.595 19.405 0.895 35.315 0.895 35.315 4.12 35.085 4.12 35.085 3.365 33.73 3.365 33.7 3.365 32.975 3.365 32.975 4.12 32.745 4.12 32.745 3.365 30.735 3.365 30.735 4.12 30.505 4.12 30.505 3.365 28.495 3.365 28.495 4.12 28.265 4.12 28.265 3.365 26.255 3.365 26.255 4.12 26.025 4.12 26.025 3.365 24.015 3.365 24.015 4.12 23.785 4.12 23.785 3.365 21.775 3.365 21.775 4.12 21.545 4.12 21.545 3.365 19.635 3.365 19.635 4.12 19.405 4.12  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.905 4.59 1.905 3.31 2.135 3.31 2.135 4.59 4.665 4.59 4.665 4.35 4.895 4.35 4.895 4.59 6.805 4.59 6.805 4.35 7.035 4.35 7.035 4.59 9.045 4.59 9.045 3.31 9.275 3.31 9.275 4.59 11.285 4.59 11.285 3.31 11.515 3.31 11.515 4.59 13.525 4.59 13.525 3.31 13.755 3.31 13.755 4.59 15.765 4.59 15.765 3.31 15.995 3.31 15.995 4.59 18.185 4.59 18.185 3.88 18.415 3.88 18.415 4.59 20.425 4.59 20.425 3.745 20.655 3.745 20.655 4.59 22.665 4.59 22.665 3.745 22.895 3.745 22.895 4.59 24.905 4.59 24.905 3.745 25.135 3.745 25.135 4.59 27.145 4.59 27.145 3.745 27.375 3.745 27.375 4.59 29.385 4.59 29.385 3.745 29.615 3.745 29.615 4.59 31.625 4.59 31.625 3.745 31.855 3.745 31.855 4.59 33.7 4.59 33.73 4.59 33.865 4.59 33.865 3.745 34.095 3.745 34.095 4.59 36.105 4.59 36.105 3.31 36.335 3.31 36.335 4.59 36.96 4.59 36.96 5.49 33.73 5.49 33.7 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 36.96 -0.45 36.96 0.45 36.435 0.45 36.435 1.49 36.205 1.49 36.205 0.45 34.25 0.45 34.25 0.665 33.91 0.665 33.91 0.45 32.01 0.45 32.01 0.665 31.67 0.665 31.67 0.45 29.77 0.45 29.77 0.665 29.43 0.665 29.43 0.45 27.53 0.45 27.53 0.665 27.19 0.665 27.19 0.45 25.29 0.45 25.29 0.665 24.95 0.665 24.95 0.45 23.05 0.45 23.05 0.665 22.71 0.665 22.71 0.45 20.81 0.45 20.81 0.665 20.47 0.665 20.47 0.45 18.515 0.45 18.515 1.49 18.285 1.49 18.285 0.45 16.095 0.45 16.095 1.49 15.865 1.49 15.865 0.45 13.855 0.45 13.855 1.49 13.625 1.49 13.625 0.45 11.615 0.45 11.615 1.455 11.385 1.455 11.385 0.45 9.43 0.45 9.43 0.64 9.09 0.64 9.09 0.45 7.19 0.45 7.19 0.64 6.85 0.64 6.85 0.45 4.95 0.45 4.95 0.64 4.61 0.64 4.61 0.45 1.595 0.45 1.595 1.16 1.365 1.16 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.885 2.505 1.805 2.505 1.805 1.62 0.245 1.62 0.245 0.68 0.475 0.68 0.475 1.39 2.035 1.39 2.035 2.505 3.65 2.505 3.65 2.735 1.115 2.735 1.115 4.12 0.885 4.12  ;
        POLYGON 5.73 3.31 8.08 3.31 8.08 1.6 5.73 1.6 5.73 1.37 8.31 1.37 8.31 2.305 16.45 2.305 16.45 2.62 8.31 2.62 8.31 3.65 5.73 3.65  ;
        POLYGON 2.925 3.31 3.155 3.31 3.155 3.89 4.405 3.89 4.405 1.595 3.55 1.595 3.55 1.365 4.635 1.365 4.635 3.89 8.585 3.89 8.585 2.85 17.065 2.85 17.065 2.505 33.7 2.505 33.7 2.735 17.295 2.735 17.295 4.12 17.065 4.12 17.065 3.08 14.875 3.08 14.875 4.12 14.645 4.12 14.645 3.08 12.635 3.08 12.635 4.12 12.405 4.12 12.405 3.08 10.395 3.08 10.395 4.12 10.165 4.12 10.165 3.08 8.815 3.08 8.815 4.12 2.925 4.12  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.905 10.265 0.905 10.265 0.68 10.5 0.68 10.5 1.75 12.505 1.75 12.505 0.68 12.735 0.68 12.735 1.75 14.745 1.75 14.745 0.68 14.975 0.68 14.975 1.75 17.165 1.75 17.165 0.68 17.395 0.68 17.395 1.75 18.8 1.75 18.8 1.865 33.73 1.865 33.73 2.095 18.61 2.095 18.61 2.075 10.27 2.075 10.27 1.135 3.32 1.135 3.32 1.865 4.175 1.865 4.175 3.65 3.945 3.65 3.945 2.095 3.09 2.095 3.09 1.49 2.485 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_16
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.2 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.065 1.21 4.33 1.21 4.33 2.15 4.065 2.15  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.575 1.015 1.575 1.015 2.71 0.71 2.71  ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.605 0.68 9.93 0.68 9.93 4.08 9.605 4.08  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.27 1.595 3.27 1.595 4.59 2.315 4.59 3.485 4.59 3.485 3.27 3.715 3.27 3.715 4.59 7.465 4.59 7.465 3.27 7.695 3.27 7.695 4.59 9.115 4.59 10.625 4.59 10.625 3.27 10.855 3.27 10.855 4.59 11.2 4.59 11.2 5.49 9.115 5.49 2.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.2 -0.45 11.2 0.45 10.955 0.45 10.955 1.49 10.725 1.49 10.725 0.45 7.995 0.45 7.995 0.885 7.765 0.885 7.765 0.45 3.615 0.45 3.615 1.02 3.385 1.02 3.385 0.45 1.595 0.45 1.595 0.895 1.365 0.895 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.115 1.155 1.115 1.155 1.125 2.315 1.125 2.315 1.915 2.085 1.915 2.085 1.355 1.085 1.355 1.085 1.345 0.475 1.345 0.475 3.27 0.575 3.27 0.575 4.08 0.245 4.08  ;
        POLYGON 2.665 0.68 2.895 0.68 2.895 2.38 4.665 2.38 4.665 1.575 4.895 1.575 4.895 2.38 5.755 2.38 5.755 2.95 5.525 2.95 5.525 2.61 2.895 2.61 2.895 4.08 2.665 4.08  ;
        POLYGON 5.245 3.18 5.985 3.18 5.985 1.225 5.345 1.225 5.345 0.885 6.19 0.885 6.19 1.115 8.435 1.115 8.435 1.915 8.205 1.915 8.205 1.345 6.215 1.345 6.215 3.41 5.475 3.41 5.475 4.08 5.245 4.08  ;
        POLYGON 7.085 1.575 7.315 1.575 7.315 2.145 8.665 2.145 8.665 0.975 9.115 0.975 9.115 2.365 8.735 2.365 8.735 4.08 8.485 4.08 8.485 2.375 7.085 2.375  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.065 1.21 4.33 1.21 4.33 2.15 4.065 2.15  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.575 1.015 1.575 1.015 2.71 0.71 2.71  ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.23 1.21 10.725 1.21 10.725 0.68 11.05 0.68 11.05 4.235 10.675 4.235 10.675 1.59 10.23 1.59  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.315 4.59 3.485 4.59 3.485 3.425 3.715 3.425 3.715 4.59 7.465 4.59 7.465 3.425 7.695 3.425 7.695 4.59 9.115 4.59 9.655 4.59 9.655 3.425 9.885 3.425 9.885 4.59 11.695 4.59 11.695 3.425 11.925 3.425 11.925 4.59 12.32 4.59 12.32 5.49 9.115 5.49 2.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 12.075 0.45 12.075 1.49 11.845 1.49 11.845 0.45 9.835 0.45 9.835 1.49 9.605 1.49 9.605 0.45 7.995 0.45 7.995 0.885 7.765 0.885 7.765 0.45 3.615 0.45 3.615 1.02 3.385 1.02 3.385 0.45 1.595 0.45 1.595 0.895 1.365 0.895 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.115 1.155 1.115 1.155 1.125 2.315 1.125 2.315 1.915 2.085 1.915 2.085 1.355 1.085 1.355 1.085 1.345 0.475 1.345 0.475 3.425 0.575 3.425 0.575 4.235 0.245 4.235  ;
        POLYGON 2.665 0.68 2.895 0.68 2.895 2.38 4.665 2.38 4.665 1.575 4.895 1.575 4.895 2.38 5.755 2.38 5.755 2.95 5.525 2.95 5.525 2.61 2.895 2.61 2.895 4.235 2.665 4.235  ;
        POLYGON 5.245 3.18 5.985 3.18 5.985 1.315 5.345 1.315 5.345 0.975 6.1 0.975 6.1 1.115 8.435 1.115 8.435 1.915 8.205 1.915 8.205 1.345 6.215 1.345 6.215 3.41 5.475 3.41 5.475 4.235 5.245 4.235  ;
        POLYGON 7.085 1.575 7.315 1.575 7.315 2.145 8.665 2.145 8.665 0.975 9.115 0.975 9.115 2.365 8.735 2.365 8.735 4.235 8.485 4.235 8.485 2.375 7.085 2.375  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.21 4.33 1.21 4.33 2.15 4.07 2.15  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.02 1.77 1.02 2.71 0.71 2.71  ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.01 1.92 11.31 1.92 11.31 0.68 11.54 0.68 11.54 1.21 13.55 1.21 13.55 0.68 13.78 0.68 13.78 1.49 13.28 1.49 13.28 4.065 13.05 4.065 13.05 1.44 11.61 1.44 11.61 2.15 11.24 2.15 11.24 4.065 11.01 4.065  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.37 4.59 1.37 3.255 1.6 3.255 1.6 4.59 2.22 4.59 3.79 4.59 3.79 3.255 4.02 3.255 4.02 4.59 7.77 4.59 7.77 3.255 8 3.255 8 4.59 9.12 4.59 9.81 4.59 9.81 3.255 10.04 3.255 10.04 4.59 12.03 4.59 12.03 3.255 12.26 3.255 12.26 4.59 14.07 4.59 14.07 3.255 14.3 3.255 14.3 4.59 15.68 4.59 15.68 5.49 9.12 5.49 2.22 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 14.9 0.45 14.9 1.49 14.67 1.49 14.67 0.45 12.66 0.45 12.66 0.98 12.43 0.98 12.43 0.45 10.24 0.45 10.24 1.02 10.01 1.02 10.01 0.45 8 0.45 8 1.02 7.77 1.02 7.77 0.45 3.62 0.45 3.62 1.02 3.39 1.02 3.39 0.45 1.6 0.45 1.6 1.02 1.37 1.02 1.37 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 0.68 0.48 0.68 0.48 1.31 2.22 1.31 2.22 2.15 1.99 2.15 1.99 1.54 0.48 1.54 0.48 3.255 0.58 3.255 0.58 4.065 0.25 4.065  ;
        POLYGON 2.57 0.68 2.9 0.68 2.9 2.38 4.67 2.38 4.67 1.81 4.9 1.81 4.9 2.38 6.06 2.38 6.06 2.72 2.8 2.72 2.8 4.065 2.57 4.065  ;
        POLYGON 5.55 2.95 6.29 2.95 6.29 1.02 5.35 1.02 5.35 0.68 7.54 0.68 7.54 1.25 8.44 1.25 8.44 2.15 8.21 2.15 8.21 1.48 7.31 1.48 7.31 0.91 6.52 0.91 6.52 3.18 5.78 3.18 5.78 4.065 5.55 4.065  ;
        POLYGON 7.33 1.81 7.56 1.81 7.56 2.38 8.89 2.38 8.89 0.68 9.12 0.68 9.12 4.065 8.79 4.065 8.79 2.61 7.33 2.61  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.88 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.295 1.77 3.295 2.71 2.95 2.71  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.21 0.97 1.21 0.97 1.31 3.905 1.31 3.905 1.495 5.195 1.495 5.195 2.44 5.5 2.44 5.5 2.67 4.965 2.67 4.965 1.725 4.135 1.725 4.135 2.295 3.675 2.295 3.675 1.54 0.97 1.54 0.97 2.295 0.705 2.295  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.455 1.77 2.455 2.71 1.83 2.71  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.91 0.845 12.355 0.845 12.355 4.36 11.91 4.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.55 1.495 3.55 1.495 4.59 3.025 4.59 3.025 3.86 3.255 3.86 3.255 4.59 6.63 4.59 6.63 3.55 6.86 3.55 6.86 4.59 9.215 4.59 9.215 3.55 9.445 3.55 9.445 4.59 9.835 4.59 11.055 4.59 11.055 3.875 11.285 3.875 11.285 4.59 11.62 4.59 12.88 4.59 12.88 5.49 11.62 5.49 9.835 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.88 -0.45 12.88 0.45 11.235 0.45 11.235 1.605 11.005 1.605 11.005 0.45 9.395 0.45 9.395 1.135 9.165 1.135 9.165 0.45 7.375 0.45 7.375 1.135 7.145 1.135 7.145 0.45 1.65 0.45 1.65 1.08 1.31 1.08 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.795 0.475 0.795 0.475 2.94 4.505 2.94 4.505 1.955 4.735 1.955 4.735 3.17 0.475 3.17 0.475 4.36 0.245 4.36  ;
        POLYGON 2.005 3.4 5.015 3.4 5.015 4.13 5.73 4.13 5.73 1.495 6.45 1.495 6.45 1.135 4.345 1.135 4.345 0.795 6.68 0.795 6.68 1.535 7.78 1.535 7.78 2.295 7.55 2.295 7.55 1.765 6.55 1.765 6.55 1.725 5.96 1.725 5.96 4.36 4.785 4.36 4.785 3.63 2.235 3.63 2.235 4.36 2.005 4.36  ;
        POLYGON 6.19 1.955 6.42 1.955 6.42 2.525 8.01 2.525 8.01 2.065 8.445 2.065 8.445 0.795 8.675 0.795 8.675 1.955 9.835 1.955 9.835 2.295 8.24 2.295 8.24 4.36 7.83 4.36 7.83 2.755 6.19 2.755  ;
        POLYGON 10.235 1.225 10.515 1.225 10.515 2.03 11.62 2.03 11.62 2.26 10.465 2.26 10.465 4.36 10.235 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.26 1.77 3.26 2.71 2.95 2.71  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.895 1.835 1.37 1.835 1.37 1.31 4.07 1.31 4.07 1.21 4.33 1.21 4.33 1.78 5 1.78 5 2.765 5.38 2.765 5.38 2.995 4.77 2.995 4.77 2.15 4.07 2.15 4.07 1.54 1.6 1.54 1.6 2.065 0.895 2.065  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.475 1.77 2.475 2.065 2.09 2.065 2.09 2.71 1.83 2.71  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.355 0.845 12.73 0.845 12.73 4.36 12.355 4.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.39 4.59 1.39 3.55 1.62 3.55 1.62 4.59 3.13 4.59 3.13 3.86 3.36 3.86 3.36 4.59 6.65 4.59 6.65 3.69 6.88 3.69 6.88 4.59 9.42 4.59 9.42 3.55 9.65 3.55 9.65 4.59 10.04 4.59 11.335 4.59 11.335 3.88 11.565 3.88 11.565 4.59 12.01 4.59 13.375 4.59 13.375 3.88 13.605 3.88 13.605 4.59 14 4.59 14 5.49 12.01 5.49 10.04 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14 -0.45 14 0.45 13.755 0.45 13.755 1.605 13.525 1.605 13.525 0.45 11.515 0.45 11.515 1.605 11.285 1.605 11.285 0.45 9.6 0.45 9.6 1.135 9.37 1.135 9.37 0.45 7.58 0.45 7.58 1.135 7.35 1.135 7.35 0.45 1.775 0.45 1.775 1.08 1.435 1.08 1.435 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.37 0.795 0.6 0.795 0.6 2.94 4.31 2.94 4.31 2.38 4.54 2.38 4.54 3.17 0.6 3.17 0.6 4.36 0.37 4.36  ;
        POLYGON 2.11 3.4 5.12 3.4 5.12 3.8 5.61 3.8 5.61 1.135 4.55 1.135 4.55 0.795 6.67 0.795 6.67 1.365 7.98 1.365 7.98 2.12 7.75 2.12 7.75 1.595 6.44 1.595 6.44 1.025 5.84 1.025 5.84 4.03 4.89 4.03 4.89 3.63 2.34 3.63 2.34 4.03 2.11 4.03  ;
        POLYGON 6.07 1.78 6.3 1.78 6.3 1.89 7.52 1.89 7.52 2.35 8.21 2.35 8.21 0.795 8.88 0.795 8.88 1.78 10.04 1.78 10.04 2.12 8.44 2.12 8.44 4.36 7.895 4.36 7.895 2.58 7.29 2.58 7.29 2.12 6.07 2.12  ;
        POLYGON 10.44 1.225 10.72 1.225 10.72 1.835 12.01 1.835 12.01 2.065 10.67 2.065 10.67 4.36 10.44 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.5 1.77 3.77 1.77 3.77 2.72 3.5 2.72  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 1.31 4.26 1.31 4.26 1.355 5.19 1.355 5.19 1.21 5.45 1.21 5.45 1.92 5.87 1.92 5.87 2.72 5.64 2.72 5.64 2.15 5.19 2.15 5.19 1.585 4.35 1.585 4.35 2.72 4.12 2.72 4.12 1.54 0.97 1.54 0.97 2.72 0.74 2.72  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.77 2.65 1.77 2.65 2.72 2.39 2.72  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.035 0.785 14.41 0.785 14.41 1.825 16.325 1.825 16.325 0.785 16.555 0.785 16.555 2.055 14.41 2.055 14.41 3.415 16.305 3.415 16.305 4.36 16.075 4.36 16.075 3.645 14.265 3.645 14.265 4.36 14.035 4.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.32 4.59 1.32 3.55 1.55 3.55 1.55 4.59 3.24 4.59 3.24 3.87 3.47 3.87 3.47 4.59 7.61 4.59 7.61 3.7 7.84 3.7 7.84 4.59 9.88 4.59 9.88 3.55 10.11 3.55 10.11 4.59 10.84 4.59 12.07 4.59 12.07 3.55 12.3 3.55 12.3 4.59 13.015 4.59 13.015 3.875 13.245 3.875 13.245 4.59 13.74 4.59 15.055 4.59 15.055 3.875 15.285 3.875 15.285 4.59 17.095 4.59 17.095 3.875 17.325 3.875 17.325 4.59 17.92 4.59 17.92 5.49 13.74 5.49 10.84 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.675 0.45 17.675 1.595 17.445 1.595 17.445 0.45 15.435 0.45 15.435 1.595 15.205 1.595 15.205 0.45 13.195 0.45 13.195 1.595 12.965 1.595 12.965 0.45 12.45 0.45 12.45 1.125 12.22 1.125 12.22 0.45 10.21 0.45 10.21 1.125 9.98 1.125 9.98 0.45 7.97 0.45 7.97 1.125 7.74 1.125 7.74 0.45 1.685 0.45 1.685 1.07 1.345 1.07 1.345 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.28 0.785 0.51 0.785 0.51 2.95 5.04 2.95 5.04 2.38 5.27 2.38 5.27 3.18 0.53 3.18 0.53 4.36 0.28 4.36  ;
        POLYGON 2.22 3.41 5.55 3.41 5.55 3.81 6.1 3.81 6.1 0.98 4.81 0.98 4.81 1.125 4.58 1.125 4.58 0.75 6.33 0.75 6.33 1.92 8.46 1.92 8.46 2.72 8.23 2.72 8.23 2.15 6.33 2.15 6.33 4.04 5.32 4.04 5.32 3.64 2.45 3.64 2.45 4.04 2.22 4.04  ;
        POLYGON 7.17 2.38 7.4 2.38 7.4 2.95 8.86 2.95 8.86 0.785 9.09 0.785 9.09 2.95 10.61 2.95 10.61 2.38 10.84 2.38 10.84 3.18 9.04 3.18 9.04 4.36 8.81 4.36 8.81 3.18 7.17 3.18  ;
        POLYGON 11.05 3.55 11.095 3.55 11.095 0.785 11.33 0.785 11.33 2.435 13.74 2.435 13.74 2.665 11.325 2.665 11.325 4.36 11.05 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 13.44 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.335 1.77 3.335 2.71 2.95 2.71  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 2.275 1.37 2.275 1.37 1.31 4.175 1.31 4.175 1.77 5.495 1.77 5.495 2.56 5.265 2.56 5.265 2.15 4.175 2.15 4.175 2.56 3.945 2.56 3.945 1.54 1.6 1.54 1.6 2.505 0.705 2.505  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.495 1.77 2.495 2.71 1.83 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.55 1.77 8.875 1.77 8.875 2.71 8.55 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.425 0.845 12.735 0.845 12.735 4.21 12.425 4.21  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.4 1.495 3.4 1.495 4.59 3.065 4.59 3.065 3.89 3.295 3.89 3.295 4.59 6.645 4.59 6.645 3.89 6.875 3.89 6.875 4.59 7.315 4.59 8.925 4.59 8.925 3.4 9.155 3.4 9.155 4.59 11.225 4.59 11.225 3.43 11.455 3.43 11.455 4.59 11.915 4.59 13.44 4.59 13.44 5.49 11.915 5.49 7.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 13.44 -0.45 13.44 0.45 11.615 0.45 11.615 1.165 11.385 1.165 11.385 0.45 7.47 0.45 7.47 1.075 7.13 1.075 7.13 0.45 1.595 0.45 1.595 1.08 1.365 1.08 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 2.94 4.545 2.94 4.545 2.38 4.775 2.38 4.775 3.17 0.475 3.17 0.475 4.21 0.245 4.21  ;
        POLYGON 2.045 3.4 7.085 3.4 7.085 3.02 5.725 3.02 5.725 1.13 4.385 1.13 4.385 0.79 5.955 0.79 5.955 2.79 7.315 2.79 7.315 3.63 5.055 3.63 5.055 4.21 4.825 4.21 4.825 3.63 2.275 3.63 2.275 4.21 2.045 4.21  ;
        POLYGON 7.905 2.94 9.325 2.94 9.325 1.54 6.415 1.54 6.415 2.56 6.185 2.56 6.185 1.31 9.325 1.31 9.325 0.79 9.555 0.79 9.555 2.22 10.715 2.22 10.715 2.56 9.555 2.56 9.555 3.17 8.135 3.17 8.135 4.21 7.905 4.21  ;
        POLYGON 10.205 2.97 11.685 2.97 11.685 1.655 10.045 1.655 10.045 1.315 10.275 1.315 10.275 1.425 11.915 1.425 11.915 3.2 10.435 3.2 10.435 4.21 10.205 4.21  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.02 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.275 3.81 2.275 3.81 2.505 3.21 2.505 3.21 3.27 2.95 3.27  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.322 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.925 1.76 6.115 1.76 6.115 2.56 5.885 2.56 5.885 1.99 4.755 1.99 4.755 2.71 4.07 2.71 4.07 1.99 1.155 1.99 1.155 2.56 0.925 2.56  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.44 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.275 2.65 2.275 2.65 2.71 1.83 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.302 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.11 1.77 9.535 1.77 9.535 2.71 9.11 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.47 1.21 12.945 1.21 12.945 0.79 13.175 0.79 13.175 4.31 12.945 4.31 12.945 2.15 12.47 2.15  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.88 1.595 3.88 1.595 4.59 3.425 4.59 3.425 4.42 3.655 4.42 3.655 4.59 7.565 4.59 7.565 3.5 7.795 3.5 7.795 4.59 8.235 4.59 9.985 4.59 9.985 3.88 10.215 3.88 10.215 4.59 11.825 4.59 11.825 3.88 12.055 3.88 12.055 4.59 12.24 4.59 14.065 4.59 14.065 3.88 14.295 3.88 14.295 4.59 14.56 4.59 14.56 5.49 12.24 5.49 8.235 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 14.295 0.45 14.295 1.6 14.065 1.6 14.065 0.45 12.055 0.45 12.055 1.53 11.825 1.53 11.825 0.45 7.835 0.45 7.835 1.13 7.605 1.13 7.605 0.45 1.815 0.45 1.815 1.13 1.585 1.13 1.585 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.695 0.79 0.695 3.42 2.665 3.42 2.665 3.5 5.125 3.5 5.125 2.22 5.355 2.22 5.355 3.73 2.49 3.73 2.49 3.65 0.475 3.65 0.475 4.31 0.245 4.31  ;
        POLYGON 2.085 3.88 2.315 3.88 2.315 3.96 5.605 3.96 5.605 2.79 6.345 2.79 6.345 1.13 4.805 1.13 4.805 0.79 6.575 0.79 6.575 2.79 8.005 2.79 8.005 2.22 8.235 2.22 8.235 3.02 5.835 3.02 5.835 4.31 5.605 4.31 5.605 4.19 2.315 4.19 2.315 4.22 2.085 4.22  ;
        POLYGON 8.865 3.42 9.765 3.42 9.765 1.54 8.21 1.54 8.21 1.99 7.365 1.99 7.365 2.56 7.135 2.56 7.135 1.76 7.98 1.76 7.98 1.31 9.745 1.31 9.745 0.79 9.995 0.79 9.995 2.22 11.375 2.22 11.375 2.56 9.995 2.56 9.995 3.65 9.095 3.65 9.095 4.31 8.865 4.31  ;
        POLYGON 10.705 3.42 12.01 3.42 12.01 1.99 10.705 1.99 10.705 0.79 10.935 0.79 10.935 1.76 12.24 1.76 12.24 3.65 10.935 3.65 10.935 4.31 10.705 4.31  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.5 1.77 3.5 2.195 3.21 2.195 3.21 2.71 2.95 2.71  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 1.965 1.83 1.965 1.83 1.31 4.285 1.31 4.285 1.89 4.755 1.89 4.755 2.875 5.37 2.875 5.37 3.105 4.525 3.105 4.525 2.12 4.055 2.12 4.055 1.54 2.09 1.54 2.09 2.71 1.83 2.71 1.83 2.195 0.97 2.195  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.375 1.77 2.65 1.77 2.65 2.71 2.375 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.55 1.77 8.985 1.77 8.985 2.71 8.55 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.265 3.42 13.515 3.42 13.515 0.845 13.745 0.845 13.745 1.92 15.27 1.92 15.27 1.21 15.755 1.21 15.755 0.845 15.985 0.845 15.985 1.655 15.53 1.655 15.53 2.15 13.745 2.15 13.745 3.42 15.535 3.42 15.535 4.29 15.305 4.29 15.305 3.65 13.495 3.65 13.495 4.29 13.265 4.29  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.305 4.59 1.305 3.48 1.535 3.48 1.535 4.59 3.045 4.59 3.045 4.12 3.275 4.12 3.275 4.59 6.565 4.59 6.565 3.48 6.795 3.48 6.795 4.59 7.535 4.59 8.785 4.59 8.785 3.65 9.015 3.65 9.015 4.59 10.205 4.59 10.205 3.88 10.435 3.88 10.435 4.59 11.065 4.59 12.245 4.59 12.245 3.88 12.475 3.88 12.475 4.59 12.915 4.59 14.285 4.59 14.285 3.88 14.515 3.88 14.515 4.59 16.325 4.59 16.325 3.88 16.555 3.88 16.555 4.59 17.36 4.59 17.36 5.49 12.915 5.49 11.065 5.49 7.535 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 17.105 0.45 17.105 1.165 16.875 1.165 16.875 0.45 14.865 0.45 14.865 1.165 14.635 1.165 14.635 0.45 12.625 0.45 12.625 1.165 12.395 1.165 12.395 0.45 10.385 0.45 10.385 1.165 10.155 1.165 10.155 0.45 7.58 0.45 7.58 1.08 7.24 1.08 7.24 0.45 1.8 0.45 1.8 1.08 1.46 1.08 1.46 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.285 0.795 0.625 0.795 0.625 2.94 4.065 2.94 4.065 2.38 4.295 2.38 4.295 3.17 0.515 3.17 0.515 4.29 0.285 4.29  ;
        POLYGON 2.025 3.48 4.82 3.48 4.82 3.335 5.6 3.335 5.6 2.655 5.535 2.655 5.535 1.135 4.495 1.135 4.495 0.795 5.765 0.795 5.765 2.49 7.305 2.49 7.305 1.935 7.535 1.935 7.535 2.72 5.83 2.72 5.83 3.565 5.035 3.565 5.035 4.29 4.805 4.29 4.805 3.71 2.255 3.71 2.255 4.29 2.025 4.29  ;
        POLYGON 7.765 3.19 9.435 3.19 9.435 1.54 6.365 1.54 6.365 2.26 6.135 2.26 6.135 1.31 9.435 1.31 9.435 0.795 9.665 0.795 9.665 1.91 11.065 1.91 11.065 2.25 9.665 2.25 9.665 3.42 7.995 3.42 7.995 4.29 7.765 4.29  ;
        POLYGON 11.225 2.53 12.685 2.53 12.685 1.655 11.275 1.655 11.275 0.845 11.505 0.845 11.505 1.425 12.915 1.425 12.915 2.76 11.455 2.76 11.455 4.29 11.225 4.29  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.21 2.27 1.21 2.27 2.16 1.83 2.16  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.015 1.77 1.015 2.39 3.065 2.39 3.065 1.83 4.03 1.83 4.03 3.2 3.69 3.2 3.69 2.09 3.295 2.09 3.295 2.62 0.71 2.62  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.87 1.21 7.21 1.21 7.21 2.16 6.87 2.16  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.72 0.845 11.05 0.845 11.05 4.23 10.72 4.23  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.42 1.595 3.42 1.595 4.59 2.955 4.59 5.225 4.59 5.225 3.42 5.455 3.42 5.455 4.59 7.685 4.59 7.685 3.42 7.915 3.42 7.915 4.59 9.57 4.59 9.57 3.42 9.8 3.42 9.8 4.59 10.37 4.59 11.76 4.59 11.76 5.49 10.37 5.49 2.955 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 9.93 0.45 9.93 1.22 9.7 1.22 9.7 0.45 5.695 0.45 5.695 1.185 5.465 1.185 5.465 0.45 1.595 0.45 1.595 1.185 1.365 1.185 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 2.85 2.955 2.85 2.955 3.19 0.575 3.19 0.575 4.23 0.245 4.23  ;
        POLYGON 3.305 3.42 3.535 3.42 3.535 4 4.26 4 4.26 1.185 3.505 1.185 3.505 0.845 5.235 0.845 5.235 1.415 6.315 1.415 6.315 2.215 6.085 2.215 6.085 1.645 5.005 1.645 5.005 1.075 4.49 1.075 4.49 4.23 3.305 4.23  ;
        POLYGON 4.785 1.875 5.855 1.875 5.855 2.445 6.745 2.445 6.745 2.39 7.605 2.39 7.605 0.845 7.835 0.845 7.835 1.875 9.025 1.875 9.025 2.215 7.835 2.215 7.835 2.62 6.895 2.62 6.895 4.23 6.665 4.23 6.665 2.675 5.625 2.675 5.625 2.215 4.785 2.215  ;
        POLYGON 8.5 2.975 9.255 2.975 9.255 1.79 9.24 1.79 9.24 1.225 8.355 1.225 8.355 0.885 9.47 0.885 9.47 1.705 10.37 1.705 10.37 2.215 10.14 2.215 10.14 1.935 9.485 1.935 9.485 3.205 8.73 3.205 8.73 4.23 8.5 4.23  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.21 2.09 1.21 2.09 2.335 1.83 2.335  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.925 1.995 1.155 1.995 1.155 2.565 2.95 2.565 2.95 1.77 3.21 1.77 3.21 2.05 3.465 2.05 3.465 3.09 4.08 3.09 4.08 3.32 3.235 3.32 3.235 2.795 0.925 2.795  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.87 1.77 7.155 1.77 7.155 2.71 6.87 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.575 0.68 11.05 0.68 11.05 2.15 10.805 2.15 10.805 4.2 10.575 4.2  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.415 4.59 1.415 3.665 1.645 3.665 1.645 4.59 3.005 4.59 5.115 4.59 5.115 3.55 5.345 3.55 5.345 4.59 7.335 4.59 7.335 3.55 7.565 3.55 7.565 4.59 9.555 4.59 9.555 3.86 9.785 3.86 9.785 4.59 10.225 4.59 11.595 4.59 11.595 3.55 11.825 3.55 11.825 4.59 12.32 4.59 12.32 5.49 10.225 5.49 3.005 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 12.075 0.45 12.075 1.49 11.845 1.49 11.845 0.45 9.835 0.45 9.835 1.305 9.605 1.305 9.605 0.45 5.695 0.45 5.695 1.02 5.465 1.02 5.465 0.45 1.595 0.45 1.595 1.02 1.365 1.02 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 3.025 3.005 3.025 3.005 3.365 0.625 3.365 0.625 4.36 0.245 4.36  ;
        POLYGON 3.355 3.55 3.585 3.55 3.585 4.13 4.31 4.13 4.31 1.765 3.505 1.765 3.505 0.68 3.735 0.68 3.735 1.535 5.965 1.535 5.965 2.335 5.735 2.335 5.735 1.765 4.54 1.765 4.54 4.36 3.355 4.36  ;
        POLYGON 5.025 1.995 5.255 1.995 5.255 2.94 8.975 2.94 8.975 2.225 7.605 2.225 7.605 0.68 7.835 0.68 7.835 1.995 9.205 1.995 9.205 3.17 6.545 3.17 6.545 4.2 6.315 4.2 6.315 3.17 5.025 3.17  ;
        POLYGON 8.535 3.4 9.995 3.4 9.995 1.765 8.485 1.765 8.485 0.68 8.715 0.68 8.715 1.535 10.225 1.535 10.225 3.63 8.765 3.63 8.765 4.21 8.535 4.21  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.245 1.21 2.65 1.21 2.65 2.15 2.245 2.15  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.945 1.92 2.015 1.92 2.015 2.38 2.88 2.38 2.88 1.92 3.22 1.92 3.22 2.33 3.77 2.33 3.77 2.945 4.195 2.945 4.195 3.27 3.51 3.27 3.51 2.61 1.785 2.61 1.785 2.15 0.945 2.15  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.87 1.77 7.23 1.77 7.23 2.71 6.87 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.51 3.09 11.76 3.09 11.76 0.84 11.99 0.84 11.99 1.21 14 1.21 14 0.84 14.23 0.84 14.23 1.65 13.85 1.65 13.85 2.15 13.59 2.15 13.59 1.44 11.99 1.44 11.99 3.09 13.78 3.09 13.78 4.25 13.55 4.25 13.55 3.32 11.74 3.32 11.74 4.25 11.51 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.61 4.59 1.61 3.705 1.84 3.705 1.84 4.59 3.28 4.59 5.39 4.59 5.39 3.55 5.62 3.55 5.62 4.59 7.61 4.59 7.61 3.875 7.84 3.875 7.84 4.59 8.45 4.59 8.45 3.875 8.68 3.875 8.68 4.59 9.07 4.59 10.49 4.59 10.49 3.875 10.72 3.875 10.72 4.59 11.3 4.59 12.53 4.59 12.53 3.55 12.76 3.55 12.76 4.59 14.57 4.59 14.57 3.875 14.8 3.875 14.8 4.59 15.68 4.59 15.68 5.49 11.3 5.49 9.07 5.49 3.28 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 15.35 0.45 15.35 1.16 15.12 1.16 15.12 0.45 13.11 0.45 13.11 0.69 12.88 0.69 12.88 0.45 10.87 0.45 10.87 1.16 10.64 1.16 10.64 0.45 8.63 0.45 8.63 1.16 8.4 1.16 8.4 0.45 5.77 0.45 5.77 1.31 5.54 1.31 5.54 0.45 1.67 0.45 1.67 1.305 1.44 1.305 1.44 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.32 0.88 0.55 0.88 0.55 2.66 0.815 2.66 0.815 2.84 3.28 2.84 3.28 3.18 0.82 3.18 0.82 4.36 0.59 4.36 0.59 2.89 0.32 2.89  ;
        POLYGON 3.63 3.55 3.86 3.55 3.86 4.13 4.425 4.13 4.425 1.77 3.58 1.77 3.58 0.97 3.81 0.97 3.81 1.54 6.23 1.54 6.23 2.31 6 2.31 6 1.77 4.655 1.77 4.655 4.36 3.63 4.36  ;
        POLYGON 5.1 2 5.33 2 5.33 2.905 6.715 2.905 6.715 2.94 8.84 2.94 8.84 1.65 7.68 1.65 7.68 0.84 7.91 0.84 7.91 1.42 9.07 1.42 9.07 3.17 6.82 3.17 6.82 4.25 6.59 4.25 6.59 3.135 5.1 3.135  ;
        POLYGON 9.47 0.84 9.75 0.84 9.75 1.94 11.3 1.94 11.3 2.28 9.7 2.28 9.7 4.25 9.47 4.25  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.77 5.45 1.77 5.45 2.15 4.63 2.15  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.77 2.65 1.77 2.65 2.71 2.39 2.71  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.225 1.38 3.455 1.38 3.455 2.475 5.75 2.475 5.75 1.77 6.035 1.77 6.035 3.27 5.75 3.27 5.75 2.705 3.225 2.705  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 0.72 0.575 0.72 0.575 4.235 0.15 4.235  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 2.97 1.595 2.97 1.595 4.59 3.835 4.59 5.31 4.59 5.31 3.48 5.65 3.48 5.65 4.59 6.815 4.59 7.28 4.59 7.28 5.49 6.815 5.49 3.835 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 5.695 0.45 5.695 0.99 5.465 0.99 5.465 0.45 1.595 0.45 1.595 1.06 1.365 1.06 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.16 3.545 3.605 3.545 3.605 2.965 3.835 2.965 3.835 3.775 1.93 3.775 1.93 2.055 0.87 2.055 0.87 1.825 1.93 1.825 1.93 0.775 3.79 0.775 3.79 1.005 2.16 1.005  ;
        POLYGON 3.945 1.31 6.585 1.31 6.585 0.72 6.815 0.72 6.815 3.775 6.385 3.775 6.385 1.54 4.175 1.54 4.175 2.11 3.945 2.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.4 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 1.77 6.57 1.77 6.57 2.15 5.75 2.15  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.255 1.77 3.255 2.71 2.95 2.71  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.005 1.775 4.235 1.775 4.235 2.47 6.87 2.47 6.87 1.77 7.315 1.77 7.315 2.71 4.005 2.71  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 0.68 1.595 0.68 1.595 4.36 1.27 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 5.115 4.59 6.645 4.59 6.645 3.55 6.875 3.55 6.875 4.59 7.995 4.59 8.4 4.59 8.4 5.49 7.995 5.49 5.115 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.4 -0.45 8.4 0.45 6.875 0.45 6.875 1.02 6.645 1.02 6.645 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.175 2.94 5.115 2.94 5.115 4.36 4.885 4.36 4.885 3.17 1.945 3.17 1.945 1.31 4.445 1.31 4.445 0.68 4.675 0.68 4.675 1.54 2.175 1.54  ;
        POLYGON 4.83 1.83 5.29 1.83 5.29 1.31 7.765 1.31 7.765 0.68 7.995 0.68 7.995 4.36 7.665 4.36 7.665 1.54 5.52 1.54 5.52 2.06 4.83 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.64 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.99 1.21 8.25 1.21 8.25 1.83 8.645 1.83 8.645 2.15 7.99 2.15  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.77 6.01 1.77 6.01 2.15 5.13 2.15  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.3 1.775 6.53 1.775 6.53 2.47 9.05 2.47 9.05 1.83 9.665 1.83 9.665 2.06 9.43 2.06 9.43 2.7 6.3 2.7  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5505 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.42 0.68 1.65 0.68 1.65 2.33 3.66 2.33 3.66 0.68 3.89 0.68 3.89 4.36 3.61 4.36 3.61 2.71 1.65 2.71 1.65 4.36 1.42 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.35 4.59 0.35 3.55 0.58 3.55 0.58 4.59 2.49 4.59 2.49 3.55 2.72 3.55 2.72 4.59 4.68 4.59 4.68 3.55 4.91 3.55 4.91 4.59 7.41 4.59 8.94 4.59 8.94 3.55 9.17 3.55 9.17 4.59 10.29 4.59 10.64 4.59 10.64 5.49 10.29 5.49 7.41 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.64 -0.45 10.64 0.45 9.17 0.45 9.17 1.02 8.94 1.02 8.94 0.45 5.01 0.45 5.01 1.02 4.78 1.02 4.78 0.45 2.77 0.45 2.77 1.49 2.54 1.49 2.54 0.45 0.53 0.45 0.53 1.49 0.3 1.49 0.3 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.9 2.93 7.41 2.93 7.41 4.36 7.18 4.36 7.18 3.16 4.67 3.16 4.67 2.115 4.24 2.115 4.24 1.775 4.67 1.775 4.67 1.31 6.74 1.31 6.74 0.68 6.97 0.68 6.97 1.54 4.9 1.54  ;
        POLYGON 7.125 1.83 7.53 1.83 7.53 0.75 8.71 0.75 8.71 1.25 10.06 1.25 10.06 0.68 10.29 0.68 10.29 4.36 9.96 4.36 9.96 1.48 8.48 1.48 8.48 0.98 7.76 0.98 7.76 2.06 7.125 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 1.21 14.97 1.21 14.97 2.555 14.71 2.555  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.35 1.77 11.61 1.77 11.61 2.71 11.35 2.71  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.375 1.77 4.375 2.71 4.07 2.71  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.67 3.21 1.67 3.21 1.9 2.65 1.9 2.65 2.995 2.39 2.995  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.675 1.77 8.105 1.77 8.81 1.77 8.81 3.195 8.405 3.195 8.405 2.155 8.105 2.155 7.675 2.155  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0032 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 2.33 6.025 2.33 6.025 1.59 5.75 1.59 5.75 1.21 6.255 1.21 6.255 3.175 5.75 3.175  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.44 0.525 3.44 0.525 4.59 1.595 4.59 4.725 4.59 4.725 3.865 4.955 3.865 4.955 4.59 7.035 4.59 8.105 4.59 10.935 4.59 10.935 3.44 11.165 3.44 11.165 4.59 13.305 4.59 15.015 4.59 15.015 3.44 15.245 3.44 15.245 4.59 16.665 4.59 17.36 4.59 17.36 5.49 16.665 5.49 13.305 5.49 8.105 5.49 7.035 5.49 1.595 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 15.545 0.45 15.545 1.43 15.315 1.43 15.315 0.45 11.065 0.45 11.065 1.43 10.835 1.43 10.835 0.45 4.955 0.45 4.955 1.43 4.725 1.43 4.725 0.45 0.475 0.45 0.475 1.43 0.245 1.43 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 1.09 1.595 1.09 1.595 4.17 1.365 4.17  ;
        POLYGON 3.605 1.09 3.835 1.09 3.835 3.355 3.915 3.355 3.915 3.695 3.605 3.695  ;
        POLYGON 2.16 3.225 2.895 3.225 2.895 3.94 4.265 3.94 4.265 3.405 6.755 3.405 6.755 1.155 6.985 1.155 6.985 3.36 7.035 3.36 7.035 4.17 6.805 4.17 6.805 3.635 4.495 3.635 4.495 4.17 2.665 4.17 2.665 3.455 1.93 3.455 1.93 1.145 2.77 1.145 2.77 1.375 2.16 1.375  ;
        POLYGON 5.29 0.695 8.105 0.695 8.105 1.345 7.875 1.345 7.875 0.925 7.445 0.925 7.445 2.385 8.055 2.385 8.055 4.17 7.825 4.17 7.825 2.615 7.215 2.615 7.215 0.925 5.52 0.925 5.52 1.79 5.575 1.79 5.575 2.13 5.29 2.13  ;
        POLYGON 9.5 1.09 10.145 1.09 10.145 3.695 9.915 3.695 9.915 2.315 9.5 2.315  ;
        POLYGON 11.955 1.09 12.185 1.09 12.185 3.695 11.955 3.695  ;
        POLYGON 8.845 3.425 9.04 3.425 9.04 1.43 8.995 1.43 8.995 1.09 9.27 1.09 9.27 4.005 10.475 4.005 10.475 2.98 11.625 2.98 11.625 3.94 12.975 3.94 12.975 1.09 13.305 1.09 13.305 4.17 11.395 4.17 11.395 3.21 10.705 3.21 10.705 4.235 8.845 4.235  ;
        POLYGON 13.675 1.145 14.48 1.145 14.48 1.375 13.905 1.375 13.905 3.245 14.225 3.245 14.225 4.25 13.995 4.25 13.995 3.475 13.675 3.475  ;
        POLYGON 14.135 2.215 14.365 2.215 14.365 2.785 16.435 2.785 16.435 1.09 16.665 1.09 16.665 3.015 16.265 3.015 16.265 4.17 16.035 4.17 16.035 3.015 14.135 3.015  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.95 1.21 17.21 1.21 17.21 2.03 16.95 2.03  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.59 1.77 13.85 1.77 13.85 2.39 13.59 2.39  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.05 1.015 2.05 1.015 3.27 0.71 3.27  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.625 2.05 4.89 2.05 4.89 2.71 4.625 2.71  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.36 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 1.77 3.815 1.77 3.815 2.26 3.51 2.26 3.51 2 2.515 2 2.515 2.39 2.285 2.39  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.24 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.56 1.69 9.79 1.69 9.79 1.77 10.23 1.77 10.83 1.77 10.83 2.83 10.6 2.83 10.6 2.15 10.23 2.15 9.56 2.15  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0816 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 1.2 6.755 1.2 6.755 3.38 6.31 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.25 4.59 0.25 3.08 0.48 3.08 0.48 4.59 1.595 4.59 5.285 4.59 5.285 4.07 5.515 4.07 5.515 4.59 7.545 4.59 7.545 3.08 7.775 3.08 7.775 4.59 9.005 4.59 10.23 4.59 13 4.59 13 3.08 13.23 3.08 13.23 4.59 15.43 4.59 17.34 4.59 17.34 3.08 17.57 3.08 17.57 4.59 18.79 4.59 19.04 4.59 19.04 5.49 18.79 5.49 15.43 5.49 10.23 5.49 9.005 5.49 1.595 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 17.67 0.45 17.67 1.54 17.44 1.54 17.44 0.45 13.19 0.45 13.19 1.54 12.96 1.54 12.96 0.45 7.875 0.45 7.875 1.54 7.645 1.54 7.645 0.45 5.635 0.45 5.635 1.54 5.405 1.54 5.405 0.45 0.475 0.45 0.475 1.54 0.245 1.54 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 1.2 1.595 1.2 1.595 3.89 1.365 3.89  ;
        POLYGON 4.045 1.615 4.285 1.615 4.285 1.2 4.515 1.2 4.515 1.845 4.275 1.845 4.275 3.38 4.045 3.38  ;
        POLYGON 2.055 3.61 2.725 3.61 2.725 3.08 2.955 3.08 2.955 3.61 7.085 3.61 7.085 2.62 8.64 2.62 8.64 1.21 8.87 1.21 8.87 3.08 9.005 3.08 9.005 3.89 8.64 3.89 8.64 2.85 7.315 2.85 7.315 3.84 2.955 3.84 2.955 3.89 1.825 3.89 1.825 1.255 3.45 1.255 3.45 1.485 2.055 1.485  ;
        POLYGON 7.105 1.77 8.18 1.77 8.18 0.75 10.23 0.75 10.23 1.54 10 1.54 10 0.98 9.33 0.98 9.33 2.36 9.465 2.36 9.465 3.66 9.95 3.66 9.95 3.08 10.18 3.08 10.18 3.89 9.235 3.89 9.235 2.57 9.1 2.57 9.1 0.98 8.41 0.98 8.41 2 7.335 2 7.335 2.39 7.105 2.39  ;
        POLYGON 11.68 1.2 12.21 1.2 12.21 3.89 11.68 3.89  ;
        POLYGON 14.08 1.2 14.31 1.2 14.31 3.89 14.08 3.89  ;
        POLYGON 11.12 1.2 11.41 1.2 11.41 4.12 12.54 4.12 12.54 2.62 13.69 2.62 13.69 4.12 15.17 4.12 15.17 1.2 15.43 1.2 15.43 4.35 13.46 4.35 13.46 2.85 12.77 2.85 12.77 4.35 11.12 4.35  ;
        POLYGON 15.7 1.255 16.605 1.255 16.605 1.485 15.93 1.485 15.93 2.665 16.42 2.665 16.42 3.89 16.19 3.89 16.19 2.895 15.7 2.895  ;
        POLYGON 16.16 2.05 16.72 2.05 16.72 2.26 18.56 2.26 18.56 1.2 18.79 1.2 18.79 3.89 18.46 3.89 18.46 2.49 16.57 2.49 16.57 2.435 16.16 2.435  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.19 1.21 19.45 1.21 19.45 2.03 19.19 2.03  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.83 2.15 16.09 2.15 16.09 2.71 15.83 2.71  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.7 2.33 1.08 2.33 1.08 2.71 0.7 2.71  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 2.15 4.89 2.15 4.89 2.71 4.63 2.71  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.36 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 1.77 3.885 1.77 3.885 2.22 2.58 2.22 2.58 2.71 2.35 2.71  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.24 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.79 1.945 12.47 1.945 12.47 1.21 12.73 1.21 12.73 1.945 13.135 1.945 13.135 2.83 12.905 2.83 12.905 2.175 11.79 2.175  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1632 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.59 1.23 6.82 1.23 6.82 1.8 8.83 1.8 8.83 1.21 9.37 1.21 9.37 3.38 9.075 3.38 9.075 2.03 6.825 2.03 6.825 3.38 6.59 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.41 4.59 0.41 3.04 0.64 3.04 0.64 4.59 1.66 4.59 5.355 4.59 5.355 4.07 5.585 4.07 5.585 4.59 7.835 4.59 7.835 4.07 8.065 4.07 8.065 4.59 10.095 4.59 10.095 3.44 10.325 3.44 10.325 4.59 11.655 4.59 12.675 4.59 15.245 4.59 15.245 3.4 15.475 3.4 15.475 4.59 17.675 4.59 19.585 4.59 19.585 3.04 19.815 3.04 19.815 4.59 21.035 4.59 21.28 4.59 21.28 5.49 21.035 5.49 17.675 5.49 12.675 5.49 11.655 5.49 1.66 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 19.915 0.45 19.915 1.57 19.685 1.57 19.685 0.45 15.435 0.45 15.435 1.57 15.205 1.57 15.205 0.45 10.18 0.45 10.18 1.57 9.95 1.57 9.95 0.45 7.94 0.45 7.94 1.57 7.71 1.57 7.71 0.45 5.7 0.45 5.7 1.57 5.47 1.57 5.47 0.45 0.54 0.45 0.54 1.57 0.31 1.57 0.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.43 1.23 1.66 1.23 1.66 3.85 1.43 3.85  ;
        POLYGON 4.115 1.695 4.35 1.695 4.35 1.23 4.58 1.23 4.58 1.925 4.345 1.925 4.345 3.38 4.115 3.38  ;
        POLYGON 2.12 3.61 2.79 3.61 2.79 3.04 3.02 3.04 3.02 3.61 9.635 3.61 9.635 2.98 10.87 2.98 10.87 1.23 11.1 1.23 11.1 3.04 11.655 3.04 11.655 3.85 11.425 3.85 11.425 3.27 10.945 3.27 10.945 3.21 9.865 3.21 9.865 3.84 3.02 3.84 3.02 3.85 1.89 3.85 1.89 1.285 3.515 1.285 3.515 1.515 2.12 1.515  ;
        POLYGON 11.56 2.405 12.675 2.405 12.675 3.85 12.445 3.85 12.445 2.635 11.33 2.635 11.33 1 10.64 1 10.64 2.03 9.885 2.03 9.885 2.71 9.655 2.71 9.655 1.8 10.41 1.8 10.41 0.77 12.235 0.77 12.235 1.57 12.005 1.57 12.005 1 11.56 1  ;
        POLYGON 13.925 1.23 14.455 1.23 14.455 3.85 13.925 3.85  ;
        POLYGON 16.325 1.23 16.555 1.23 16.555 3.85 16.325 3.85  ;
        POLYGON 13.125 1.23 13.695 1.23 13.695 4.08 14.785 4.08 14.785 2.94 15.935 2.94 15.935 4.08 17.445 4.08 17.445 1.23 17.675 1.23 17.675 4.31 15.705 4.31 15.705 3.17 15.015 3.17 15.015 4.31 13.465 4.31 13.465 1.57 13.125 1.57  ;
        POLYGON 17.945 1.285 18.85 1.285 18.85 1.515 18.175 1.515 18.175 2.72 18.795 2.72 18.795 3.85 18.565 3.85 18.565 2.95 17.945 2.95  ;
        POLYGON 18.405 2.15 18.635 2.15 18.635 2.26 20.805 2.26 20.805 1.23 21.035 1.23 21.035 3.85 20.705 3.85 20.705 2.49 18.405 2.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.8 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.33 2.09 2.33 2.09 3.27 1.83 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.635 1.77 0.975 1.77 0.975 2.71 0.635 2.71  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4362 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 3.02 1.53 3.02 1.53 3.6 2.32 3.6 2.32 1.59 1.27 1.59 1.27 1.21 2.29 1.21 2.29 0.68 2.55 0.68 2.55 3.83 1.27 3.83  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.25 4.59 0.25 3.69 0.48 3.69 0.48 4.59 2.29 4.59 2.29 4.16 2.52 4.16 2.52 4.59 2.8 4.59 2.8 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.8 -0.45 2.8 0.45 0.48 0.45 0.48 1.165 0.25 1.165 0.25 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.685 1.83 2.715 1.83 2.715 2.305 1.685 2.305  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.21 0.97 1.21 0.97 2.94 3.015 2.94 3.015 1.83 4.03 1.83 4.03 2.1 3.245 2.1 3.245 3.17 0.71 3.17  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3972 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 3.4 3.39 3.4 3.39 3.35 4.07 3.35 4.07 2.33 4.26 2.33 4.26 1.59 2.285 1.59 2.285 0.68 2.515 0.68 2.515 1.21 4.49 1.21 4.49 3.58 3.535 3.58 3.535 4.21 3.305 4.21 3.305 3.63 1.495 3.63 1.495 4.21 1.265 4.21  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.86 0.475 3.86 0.475 4.59 2.285 4.59 2.285 3.86 2.515 3.86 2.515 4.59 4.325 4.59 4.325 3.86 4.555 3.86 4.555 4.59 5.04 4.59 5.04 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 4.555 0.45 4.555 0.695 4.325 0.695 4.325 0.45 0.475 0.45 0.475 1.165 0.245 1.165 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.67 2.47 3.01 2.47 3.01 2.95 5.73 2.95 5.73 2.47 6.07 2.47 6.07 3.21 2.67 3.21  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.77 1.83 8.11 1.83 8.11 2.15 0.77 2.15  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.8538 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 3.55 7.385 3.55 7.385 3.23 8.34 3.23 8.34 1.105 7.94 1.105 7.94 1.1 2.275 1.1 2.275 0.87 8.145 0.87 8.145 0.875 8.57 0.875 8.57 3.46 7.75 3.46 7.75 4.33 7.37 4.33 7.37 3.78 5.575 3.78 5.575 4.36 5.345 4.36 5.345 3.78 3.535 3.78 3.535 4.36 3.305 4.36 3.305 3.78 1.495 3.78 1.495 4.36 1.265 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.69 0.475 3.69 0.475 4.59 2.285 4.59 2.285 4.16 2.515 4.16 2.515 4.59 4.325 4.59 4.325 4.16 4.555 4.16 4.555 4.59 6.365 4.59 6.365 4.16 6.595 4.16 6.595 4.59 8.405 4.59 8.405 3.69 8.635 3.69 8.635 4.59 8.96 4.59 8.96 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 8.69 0.45 8.69 0.64 8.35 0.64 8.35 0.45 4.575 0.45 4.575 0.64 4.235 0.64 4.235 0.45 0.555 0.45 0.555 1.165 0.325 1.165 0.325 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 3.92 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.21 3.21 1.21 3.21 2.15 2.95 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.71 1.83 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.33 1.105 2.33 1.105 3.27 0.71 3.27  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9824 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 3.55 2.95 3.55 2.95 2.89 3.44 2.89 3.44 0.845 3.67 0.845 3.67 3.83 1.63 3.83 1.63 4.36 1.4 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.38 4.59 0.38 3.59 0.61 3.59 0.61 4.59 2.42 4.59 2.42 4.06 2.65 4.06 2.65 4.59 3.92 4.59 3.92 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 3.92 -0.45 3.92 0.45 0.61 0.45 0.61 1.165 0.38 1.165 0.38 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand3_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.865 1.21 3.21 1.21 3.21 2.15 2.865 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 2.38 4.63 2.38 4.63 1.21 4.995 1.21 4.995 2.61 1.79 2.61  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.77 1.92 1.27 1.92 1.27 1.915 1.53 1.915 1.53 2.84 5.74 2.84 5.74 2.07 6.015 2.07 6.015 3.07 1.3 3.07 1.3 2.15 0.77 2.15  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.964 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 3.3 5.575 3.3 5.575 4.11 5.345 4.11 5.345 3.53 3.535 3.53 3.535 4.11 3.305 4.11 3.305 3.53 1.495 3.53 1.495 4.11 1.265 4.11 1.265 3.53 0.15 3.53 0.15 0.865 0.87 0.865 0.87 0.75 3.59 0.75 3.59 0.98 1.07 0.98 1.07 1.095 0.41 1.095  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 4.23 0.475 4.23 0.475 4.59 2.285 4.59 2.285 3.76 2.515 3.76 2.515 4.59 4.325 4.59 4.325 3.76 4.555 3.76 4.555 4.59 6.365 4.59 6.365 3.76 6.595 3.76 6.595 4.59 7.28 4.59 7.28 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 6.595 0.45 6.595 1.16 6.365 1.16 6.365 0.45 0.67 0.45 0.67 0.635 0.33 0.635 0.33 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand3_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.3 1.77 9.93 1.77 9.93 2.27 11.23 2.27 11.23 2.5 9.3 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.75 2.215 0.98 2.215 0.98 2.73 3.51 2.73 3.51 2.27 4.13 2.27 4.13 2.73 8.125 2.73 8.125 2.215 8.355 2.215 8.355 2.96 0.75 2.96  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 1.81 4.64 1.81 4.64 2.27 6.27 2.27 6.27 2.5 4.41 2.5 4.41 2.04 1.99 2.04 1.99 2.5 1.21 2.5  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.22 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 3.19 11.965 3.19 11.965 1.515 9.825 1.515 9.825 1.14 10.055 1.14 10.055 1.285 12.01 1.285 12.01 1.14 12.79 1.14 12.79 1.53 12.195 1.53 12.195 4.36 11.965 4.36 11.965 3.42 9.955 3.42 9.955 4.36 9.725 4.36 9.725 3.42 7.915 3.42 7.915 4.36 7.685 4.36 7.685 3.42 5.775 3.42 5.775 4.36 5.545 4.36 5.545 3.42 3.635 3.42 3.635 4.36 3.405 4.36 3.405 3.42 1.495 3.42 1.495 4.36 1.265 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.65 0.475 3.65 0.475 4.59 2.285 4.59 2.285 3.875 2.515 3.875 2.515 4.59 4.425 4.59 4.425 3.65 4.655 3.65 4.655 4.59 6.565 4.59 6.565 3.65 6.795 3.65 6.795 4.59 8.705 4.59 8.705 3.65 8.935 3.65 8.935 4.59 10.845 4.59 10.845 3.65 11.075 3.65 11.075 4.59 13.085 4.59 13.085 3.65 13.315 3.65 13.315 4.59 13.415 4.59 14 4.59 14 5.49 13.415 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14 -0.45 14 0.45 6.895 0.45 6.895 1.11 6.665 1.11 6.665 0.45 2.615 0.45 2.615 1.11 2.385 1.11 2.385 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.77 0.475 0.77 0.475 1.35 2.845 1.35 2.845 0.77 4.755 0.77 4.755 1.35 8.94 1.35 8.94 0.68 13.415 0.68 13.415 1.58 13.185 1.58 13.185 0.91 11.23 0.91 11.23 1.055 10.89 1.055 10.89 0.91 9.17 0.91 9.17 1.58 4.525 1.58 4.525 1 3.075 1 3.075 1.58 0.245 1.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nand3_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.985 2.27 4.33 2.27 4.33 2.71 3.985 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.915 2.215 3.21 2.215 3.21 2.71 2.915 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.125 1.77 1.125 2.5 0.71 2.5  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.42 3.26 3.54 3.26 3.54 3.025 4.56 3.025 4.56 1.49 4.48 1.49 4.48 0.68 4.79 0.68 4.79 3.255 3.77 3.255 3.77 4.36 3.46 4.36 3.46 3.49 1.65 3.49 1.65 4.36 1.42 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.4 4.59 0.4 3.72 0.63 3.72 0.63 4.59 2.44 4.59 2.44 3.72 2.67 3.72 2.67 4.59 4.48 4.59 4.48 3.485 4.71 3.485 4.71 4.59 5.04 4.59 5.04 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 0.63 0.45 0.63 1.49 0.4 1.49 0.4 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand4_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 2.215 3.875 2.215 3.875 2.71 3.51 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.865 2.215 3.095 2.215 3.095 2.94 4.235 2.94 4.235 2.215 6.015 2.215 6.015 2.71 4.465 2.71 4.465 3.17 2.865 3.17  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.755 7.035 1.755 7.035 2.555 6.805 2.555 6.805 1.985 2.09 1.985 2.09 2.555 1.83 2.555  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 2.215 1.27 2.215 1.27 1.77 1.53 1.77 1.53 3.31 2.235 3.31 2.235 3.4 4.695 3.4 4.695 2.94 7.825 2.94 7.825 2.215 8.055 2.215 8.055 3.17 4.925 3.17 4.925 3.63 2.05 3.63 2.05 3.54 1.3 3.54 1.3 2.555 0.825 2.555  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.8096 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.475 3.77 1.865 3.77 1.865 3.86 5.065 3.86 5.065 3.815 6.365 3.815 6.365 3.4 8.635 3.4 8.635 4.36 8.405 4.36 8.405 3.63 6.595 3.63 6.595 4.045 5.205 4.045 5.205 4.09 1.68 4.09 1.68 4 0.475 4 0.475 4.36 0.15 4.36 0.15 1.755 0.81 1.755 0.81 0.68 4.555 0.68 4.555 1.49 4.325 1.49 4.325 0.91 1.04 0.91 1.04 1.985 0.475 1.985  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 4.23 1.495 4.23 1.495 4.59 3.305 4.59 3.305 4.32 3.535 4.32 3.535 4.59 5.345 4.59 5.345 4.275 5.575 4.275 5.575 4.59 7.385 4.59 7.385 3.86 7.615 3.86 7.615 4.59 8.96 4.59 8.96 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 8.635 0.45 8.635 1.49 8.405 1.49 8.405 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand4_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.67 1.755 12.595 1.755 12.595 2.27 14.23 2.27 14.23 2.5 12.365 2.5 12.365 1.985 10.15 1.985 10.15 2.5 9.67 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.93 2.27 9.27 2.27 9.27 2.73 11.35 2.73 11.35 2.215 12.135 2.215 12.135 2.73 15.705 2.73 15.705 2.215 15.935 2.215 15.935 2.96 8.93 2.96  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.27 1.05 2.27 1.05 2.73 3.745 2.73 3.745 2.215 3.975 2.215 3.975 2.73 6.3 2.73 6.3 2.27 8.11 2.27 8.11 2.5 6.53 2.5 6.53 2.96 0.71 2.96  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.755 4.435 1.755 4.435 2.27 6.07 2.27 6.07 2.5 4.205 2.5 4.205 1.985 2.17 1.985 2.17 2.5 1.83 2.5  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.6976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 3.19 16.165 3.19 16.165 1.425 10.39 1.425 10.39 1.195 16.395 1.195 16.395 3.42 15.775 3.42 15.775 4.36 15.545 4.36 15.545 3.42 13.735 3.42 13.735 4.36 13.505 4.36 13.505 3.42 11.695 3.42 11.695 4.36 11.465 4.36 11.465 3.42 9.655 3.42 9.655 4.36 9.425 4.36 9.425 3.42 7.615 3.42 7.615 4.36 7.385 4.36 7.385 3.42 5.575 3.42 5.575 4.36 5.345 4.36 5.345 3.42 3.535 3.42 3.535 4.36 2.89 4.36 2.89 3.42 1.495 3.42 1.495 4.36 1.265 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.65 0.475 3.65 0.475 4.59 2.285 4.59 2.285 3.65 2.515 3.65 2.515 4.59 4.325 4.59 4.325 3.65 4.555 3.65 4.555 4.59 6.365 4.59 6.365 3.65 6.595 3.65 6.595 4.59 8.405 4.59 8.405 3.65 8.635 3.65 8.635 4.59 10.445 4.59 10.445 3.65 10.675 3.65 10.675 4.59 12.485 4.59 12.485 3.65 12.715 3.65 12.715 4.59 14.525 4.59 14.525 3.65 14.755 3.65 14.755 4.59 16.565 4.59 16.565 3.65 16.795 3.65 16.795 4.59 16.85 4.59 17.36 4.59 17.36 5.49 16.85 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 6.595 0.45 6.595 1.02 6.365 1.02 6.365 0.45 2.515 0.45 2.515 1.02 2.285 1.02 2.285 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.26 4.325 1.26 4.325 0.68 4.555 0.68 4.555 1.26 9.93 1.26 9.93 0.735 16.85 0.735 16.85 0.965 10.16 0.965 10.16 1.49 0.245 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nand4_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 3.36 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.68 2.27 1.02 2.27 1.02 2.71 0.68 2.71  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2836 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 0.68 1.595 0.68 1.595 2.785 2.665 2.785 2.665 4.36 2.435 4.36 2.435 3.015 1.27 3.015  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 3.36 4.59 3.36 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 3.36 -0.45 3.36 0.45 2.715 0.45 2.715 1.4 2.485 1.4 2.485 0.45 0.475 0.45 0.475 1.4 0.245 1.4 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.875 2.215 1.105 2.215 1.105 2.94 3.51 2.94 3.51 1.77 3.77 1.77 3.77 2.27 3.95 2.27 3.95 3.17 0.875 3.17  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9999 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.485 3.55 4.18 3.55 4.18 1.72 4.07 1.72 4.07 1.49 1.365 1.49 1.365 0.68 1.595 0.68 1.595 1.16 3.605 1.16 3.605 0.68 3.835 0.68 3.835 1.21 4.41 1.21 4.41 3.78 2.715 3.78 2.715 4.36 2.485 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 4.675 4.59 4.675 3.55 4.905 3.55 4.905 4.59 5.6 4.59 5.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.955 0.45 4.955 1.4 4.725 1.4 4.725 0.45 2.715 0.45 2.715 0.93 2.485 0.93 2.485 0.45 0.475 0.45 0.475 1.4 0.245 1.4 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.06 2.27 3.58 2.27 3.58 1.77 4.89 1.77 4.89 2.27 6.62 2.27 6.62 2.5 4.63 2.5 4.63 2 3.81 2 3.81 2.5 3.06 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 2.27 2.83 2.27 2.83 2.73 4.04 2.73 4.04 2.27 4.38 2.27 4.38 2.73 6.85 2.73 6.85 2.27 8.86 2.27 8.86 2.5 7.08 2.5 7.08 2.96 2.6 2.96 2.6 2.5 1.2 2.5  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.0913 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.26 1.365 1.26 1.365 0.68 1.595 0.68 1.595 1.26 3.605 1.26 3.605 0.68 3.835 0.68 3.835 1.26 5.845 1.26 5.845 0.68 6.075 0.68 6.075 1.26 8.085 1.26 8.085 0.68 8.315 0.68 8.315 1.49 0.97 1.49 0.97 3.19 7.145 3.19 7.145 4.36 6.915 4.36 6.915 3.42 2.715 3.42 2.715 4.36 2.485 4.36 2.485 3.42 0.71 3.42  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.65 0.525 3.65 0.525 4.59 4.675 4.59 4.675 3.65 4.905 3.65 4.905 4.59 9.155 4.59 9.155 3.65 9.385 3.65 9.385 4.59 10.08 4.59 10.08 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 9.435 0.45 9.435 1.4 9.205 1.4 9.205 0.45 7.195 0.45 7.195 1.02 6.965 1.02 6.965 0.45 4.955 0.45 4.955 1.02 4.725 1.02 4.725 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.21 1.77 3.21 2.555 2.95 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.5636 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.68 1.595 0.68 1.595 1.25 3.605 1.25 3.605 0.68 3.835 0.68 3.835 4.36 3.505 4.36 3.505 1.48 1.365 1.48  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 4.48 4.59 4.48 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor3_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.475 2.215 3.77 2.215 3.77 2.71 3.475 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.215 2.135 2.215 2.135 2.94 5.215 2.94 5.215 2.215 5.445 2.215 5.445 3.17 1.83 3.17  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.215 1.495 2.215 1.495 3.4 6.31 3.4 6.31 2.215 6.57 2.215 6.57 3.63 1.265 3.63  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.6514 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.21 2.485 1.21 2.485 0.68 2.715 0.68 2.715 1.25 4.725 1.25 4.725 0.68 4.955 0.68 4.955 1.25 6.965 1.25 6.965 0.68 7.195 0.68 7.195 1.48 1.035 1.48 1.035 3.93 3.84 3.93 3.84 4.16 0.805 4.16 0.805 1.59 0.245 1.59  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.875 0.575 3.875 0.575 4.59 6.865 4.59 6.865 3.875 7.095 3.875 7.095 4.59 7.84 4.59 7.84 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 6.075 0.45 6.075 1.02 5.845 1.02 5.845 0.45 3.835 0.45 3.835 1.02 3.605 1.02 3.605 0.45 1.595 0.45 1.595 0.98 1.365 0.98 1.365 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor3_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.8 1.71 11.73 1.71 11.73 2.15 9.8 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 2.325 1.055 2.325 1.055 2.895 3.51 2.895 3.51 2.33 3.77 2.33 3.77 2.38 4.33 2.38 4.33 2.895 6.745 2.895 6.745 2.38 8.81 2.38 8.81 2.61 6.975 2.61 6.975 3.125 0.825 3.125  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 1.77 6.515 1.77 6.515 2.665 6.285 2.665 6.285 2.15 4.07 2.15 4.07 2 3.28 2 3.28 2.61 2.94 2.61  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.734 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.325 2.65 11.96 2.65 11.96 1.48 1.365 1.48 1.365 0.68 1.595 0.68 1.595 1.25 3.605 1.25 3.605 0.68 3.835 0.68 3.835 1.25 5.845 1.25 5.845 0.68 6.075 0.68 6.075 1.25 8.085 1.25 8.085 0.68 8.315 0.68 8.315 1.25 10.325 1.25 10.325 0.68 10.555 0.68 10.555 1.25 12.565 1.25 12.565 0.68 12.795 0.68 12.795 1.48 12.19 1.48 12.19 3.09 12.695 3.09 12.695 3.9 11.91 3.9 11.91 2.88 10.555 2.88 10.555 3.9 10.325 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.825 2.615 3.825 2.615 4.59 6.865 4.59 6.865 3.815 7.095 3.815 7.095 4.59 13.815 4.59 14.56 4.59 14.56 5.49 13.815 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 13.915 0.45 13.915 1.02 13.685 1.02 13.685 0.45 11.675 0.45 11.675 1.02 11.445 1.02 11.445 0.45 9.435 0.45 9.435 1.02 9.205 1.02 9.205 0.45 7.195 0.45 7.195 1.02 6.965 1.02 6.965 0.45 4.955 0.45 4.955 1.02 4.725 1.02 4.725 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.11 0.475 3.11 0.475 3.355 7.605 3.355 7.605 4.13 11.345 4.13 11.345 3.11 11.575 3.11 11.575 4.13 13.585 4.13 13.585 3.11 13.815 3.11 13.815 4.36 7.375 4.36 7.375 3.585 4.855 3.585 4.855 4.165 4.625 4.165 4.625 3.585 0.475 3.585 0.475 3.92 0.245 3.92  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor3_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.555 4.07 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4916 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.68 1.595 0.68 1.595 1.21 3.605 1.21 3.605 0.68 3.835 0.68 3.835 2.785 4.855 2.785 4.855 4.36 4.625 4.36 4.625 3.015 3.51 3.015 3.51 1.44 1.365 1.44  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 5.6 4.59 5.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.955 0.45 4.955 1.005 4.725 1.005 4.725 0.45 2.715 0.45 2.715 0.98 2.485 0.98 2.485 0.45 0.475 0.45 0.475 1.005 0.245 1.005 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor4_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.87 2.15 7.13 2.15 7.13 2.71 6.87 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.77 1.77 6.57 1.77 6.57 2.94 8.89 2.94 8.89 2.215 9.12 2.215 9.12 3.17 6.34 3.17 6.34 2.555 5.77 2.555  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 2.215 1.16 2.215 1.16 2.785 4.07 2.785 4.07 1.77 4.51 1.77 4.51 3.015 0.93 3.015  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.622 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.7182 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.68 1.6 0.68 1.6 1.225 3.61 1.225 3.61 0.68 3.84 0.68 3.84 1.21 6.21 1.21 6.21 0.68 6.44 0.68 6.44 1.225 8.45 1.225 8.45 0.68 8.68 0.68 8.68 1.455 5.45 1.455 5.45 3.4 7.51 3.4 7.51 3.89 7.28 3.89 7.28 3.63 5.19 3.63 5.19 1.455 1.37 1.455  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.44 4.59 2.44 3.705 2.67 3.705 2.67 4.59 9.7 4.59 10.08 4.59 10.08 5.49 9.7 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 9.8 0.45 9.8 0.995 9.57 0.995 9.57 0.45 7.56 0.45 7.56 0.995 7.33 0.995 7.33 0.45 5.14 0.45 5.14 0.98 4.91 0.98 4.91 0.45 2.72 0.45 2.72 0.995 2.49 0.995 2.49 0.45 0.48 0.45 0.48 1.02 0.25 1.02 0.25 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.35 3.55 0.58 3.55 0.58 4.13 1.98 4.13 1.98 3.245 3.13 3.245 3.13 4.13 9.47 4.13 9.47 3.55 9.7 3.55 9.7 4.36 2.9 4.36 2.9 3.475 2.21 3.475 2.21 4.36 0.35 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor4_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.465 2.215 17.46 2.215 17.46 2.71 13.465 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.87 1.755 20.01 1.755 20.01 2.555 19.55 2.555 19.55 1.985 11.1 1.985 11.1 2.555 10.87 2.555  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.33 1.77 1.33 2.785 4.59 2.785 4.59 2.215 4.82 2.215 4.82 2.785 7.47 2.785 7.47 2.27 9.715 2.27 9.715 2.5 7.7 2.5 7.7 3.015 1.1 3.015 1.1 2.15 0.71 2.15  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.48 1.755 7.24 1.755 7.24 2.555 6.78 2.555 6.78 1.985 3.71 1.985 3.71 2.555 3.48 2.555  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.3894 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.89 3.09 20.405 3.09 20.405 1.59 20.175 1.59 20.175 1.455 6.52 1.455 6.52 0.91 5.91 0.91 5.91 1.455 1.68 1.455 1.68 0.68 1.91 0.68 1.91 1.225 3.92 1.225 3.92 0.68 4.15 0.68 4.15 1.225 5.68 1.225 5.68 0.68 6.75 0.68 6.75 1.225 8.76 1.225 8.76 0.68 8.99 0.68 8.99 1.225 11.36 1.225 11.36 0.68 11.59 0.68 11.59 1.225 13.96 1.225 13.96 0.68 14.19 0.68 14.19 1.225 16.56 1.225 16.56 0.68 16.79 0.68 16.79 1.225 19.16 1.225 19.16 0.68 19.39 0.68 19.39 1.21 20.635 1.21 20.635 3.32 18.04 3.32 18.04 3.9 17.81 3.9 17.81 3.32 13.12 3.32 13.12 3.9 12.89 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.75 4.59 2.75 3.705 2.98 3.705 2.98 4.59 7.59 4.59 7.59 3.705 7.82 3.705 7.82 4.59 20.59 4.59 21.28 4.59 21.28 5.49 20.59 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.69 0.45 20.69 0.98 20.46 0.98 20.46 0.45 18.09 0.45 18.09 0.995 17.86 0.995 17.86 0.45 15.49 0.45 15.49 0.97 15.26 0.97 15.26 0.45 12.89 0.45 12.89 0.995 12.66 0.995 12.66 0.45 10.29 0.45 10.29 0.995 10.06 0.995 10.06 0.45 7.87 0.45 7.87 0.995 7.64 0.995 7.64 0.45 5.45 0.45 5.45 0.995 5.22 0.995 5.22 0.45 3.03 0.45 3.03 0.995 2.8 0.995 2.8 0.45 0.79 0.45 0.79 0.995 0.56 0.995 0.56 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.66 3.55 0.89 3.55 0.89 4.13 2.29 4.13 2.29 3.245 8.28 3.245 8.28 4.13 15.21 4.13 15.21 3.55 15.44 3.55 15.44 4.13 20.36 4.13 20.36 3.55 20.59 3.55 20.59 4.36 8.05 4.36 8.05 3.475 5.4 3.475 5.4 4.36 5.17 4.36 5.17 3.475 2.52 3.475 2.52 4.36 0.66 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor4_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.68 2.27 1.02 2.27 1.02 2.71 0.68 2.71  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.27 3.29 2.27 3.29 2.71 2.95 2.71  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9119 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.14 1.595 1.14 1.595 2.785 2.615 2.785 2.615 4.36 2.385 4.36 2.385 3.015 1.27 3.015  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 2.715 4.59 3.585 4.59 3.585 3.55 3.815 3.55 3.815 4.59 4.48 4.59 4.48 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 3.835 0.45 3.835 1.655 3.605 1.655 3.605 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 2.715 0.68 2.715 1.655 2.485 1.655 2.485 0.91 0.475 0.91 0.475 1.655 0.245 1.655  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.035 2.215 4.33 2.215 4.33 2.71 4.035 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.27 3.31 2.27 3.31 2.94 6.285 2.94 6.285 2.215 6.515 2.215 6.515 3.17 2.95 3.17  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 2.27 1.07 2.27 1.07 2.65 0.65 2.65  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.3628 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.4 6.745 3.4 6.745 1.95 3.605 1.95 3.605 1.14 3.835 1.14 3.835 1.72 5.19 1.72 5.19 1.14 6.075 1.14 6.075 1.72 6.975 1.72 6.975 3.63 4.905 3.63 4.905 4.36 4.675 4.36 4.675 3.63 1.595 3.63 1.595 4.32 1.365 4.32  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.665 0.575 3.665 0.575 4.59 2.385 4.59 2.385 3.86 2.615 3.86 2.615 4.59 6.865 4.59 6.865 3.86 7.095 3.86 7.095 4.59 7.195 4.59 7.84 4.59 7.84 5.49 7.195 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 1.595 0.45 1.595 1.49 1.365 1.49 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.72 2.485 1.72 2.485 0.68 7.195 0.68 7.195 1.49 6.965 1.49 6.965 0.91 4.955 0.91 4.955 1.49 4.725 1.49 4.725 0.91 2.715 0.91 2.715 1.95 0.245 1.95  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.06 2.27 3.51 2.27 3.51 1.77 3.77 1.77 3.77 1.81 4.84 1.81 4.84 2.27 6.57 2.27 6.57 2.5 4.61 2.5 4.61 2.04 3.77 2.04 3.77 2.5 3.06 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.25 2.27 2.83 2.27 2.83 2.73 4.04 2.73 4.04 2.27 4.38 2.27 4.38 2.73 6.8 2.73 6.8 2.27 8.81 2.27 8.81 2.5 7.03 2.5 7.03 2.96 2.6 2.96 2.6 2.5 1.25 2.5  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.27 2.27 11.35 2.27 11.35 1.77 11.61 1.77 11.61 2.27 12.85 2.27 12.85 2.5 10.27 2.5  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.7986 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.02 3.19 12.745 3.19 12.745 4.36 12.515 4.36 12.515 3.42 10.555 3.42 10.555 4.36 10.325 4.36 10.325 3.42 7.145 3.42 7.145 4.36 6.915 4.36 6.915 3.42 2.715 3.42 2.715 4.36 2.485 4.36 2.485 3.42 0.79 3.42 0.79 1.81 1.365 1.81 1.365 1.14 1.595 1.14 1.595 1.81 2.95 1.81 2.95 1.14 4.12 1.14 4.12 1.34 5.845 1.34 5.845 1.14 6.075 1.14 6.075 1.34 8.085 1.34 8.085 1.14 8.315 1.14 8.315 1.57 3.935 1.57 3.935 1.48 3.21 1.48 3.21 2.04 1.02 2.04  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.65 0.575 3.65 0.575 4.59 4.675 4.59 4.675 3.65 4.905 3.65 4.905 4.59 9.105 4.59 9.105 3.65 9.335 3.65 9.335 4.59 11.345 4.59 11.345 3.65 11.575 3.65 11.575 4.59 13.635 4.59 13.635 3.65 13.865 3.65 13.865 4.59 13.915 4.59 14.56 4.59 14.56 5.49 13.915 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 12.795 0.45 12.795 1.11 12.565 1.11 12.565 0.45 10.555 0.45 10.555 1.195 10.325 1.195 10.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 9.435 0.68 9.435 1.425 10.95 1.425 10.95 1.31 11.445 1.31 11.445 0.73 11.905 0.73 11.905 1.35 13.685 1.35 13.685 0.77 13.915 0.77 13.915 1.58 11.775 1.58 11.775 1.54 11.15 1.54 11.15 1.655 9.205 1.655 9.205 0.91 7.195 0.91 7.195 1.11 6.965 1.11 6.965 0.91 4.955 0.91 4.955 1.11 4.725 1.11 4.725 0.91 2.715 0.91 2.715 1.58 2.485 1.58 2.485 0.91 0.475 0.91 0.475 1.58 0.245 1.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.21 1.77 3.21 2.555 2.95 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.555 4.07 2.555  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 3.27 0.71 3.27  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.535 2.785 3.51 2.785 3.51 1.14 3.835 1.14 3.835 3.015 2.765 3.015 2.765 4.36 2.535 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 4.955 4.59 5.6 4.59 5.6 5.49 4.955 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 1.595 0.45 1.595 1.525 1.365 1.525 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.715 0.475 0.715 0.475 1.755 2.485 1.755 2.485 0.68 4.955 0.68 4.955 1.525 4.725 1.525 4.725 0.91 2.715 0.91 2.715 1.985 0.245 1.985  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.28 2.27 6.62 2.27 6.62 2.71 6.28 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.35 2.27 5.69 2.27 5.69 2.94 6.87 2.94 6.87 2.215 8.755 2.215 8.755 3.17 5.35 3.17  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.75 2.27 2.09 2.27 2.09 2.71 1.75 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.27 1.21 2.27 1.21 2.94 2.39 2.94 2.39 2.27 4.33 2.27 4.33 3.17 0.87 3.17  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.7335 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.535 3.4 8.985 3.4 8.985 1.985 5.845 1.985 5.845 1.14 6.075 1.14 6.075 1.755 7.99 1.755 7.99 1.14 8.315 1.14 8.315 1.755 9.215 1.755 9.215 3.63 7.145 3.63 7.145 4.36 6.915 4.36 6.915 3.63 2.765 3.63 2.765 4.36 2.535 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.86 0.575 3.86 0.575 4.59 4.625 4.59 4.625 3.86 4.855 3.86 4.855 4.59 9.105 4.59 9.105 3.86 9.335 3.86 9.335 4.59 9.435 4.59 10.08 4.59 10.08 5.49 9.435 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 3.835 0.45 3.835 1.055 3.605 1.055 3.605 0.45 1.595 0.45 1.595 1.525 1.365 1.525 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.715 0.475 0.715 0.475 1.755 2.485 1.755 2.485 1.285 4.725 1.285 4.725 0.68 9.435 0.68 9.435 1.525 9.205 1.525 9.205 0.91 7.195 0.91 7.195 1.525 6.965 1.525 6.965 0.91 4.955 0.91 4.955 1.985 0.245 1.985  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.73 1.755 13.745 1.755 13.745 2.27 15.53 2.27 15.53 2.5 13.515 2.5 13.515 1.985 11.34 1.985 11.34 2.5 10.73 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.885 2.215 10.115 2.215 10.115 2.73 12.47 2.73 12.47 2.215 13.285 2.215 13.285 2.73 17.485 2.73 17.485 2.215 17.715 2.215 17.715 2.96 9.885 2.96  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.11 1.77 5.04 1.77 5.04 2.27 6.57 2.27 6.57 2.5 4.81 2.5 4.81 2.15 4.58 2.15 4.58 2.04 3.45 2.04 3.45 2.5 3.11 2.5  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.875 2.215 1.105 2.215 1.105 2.73 4.04 2.73 4.04 2.27 4.38 2.27 4.38 2.73 6.8 2.73 6.8 2.27 8.81 2.27 8.81 2.5 7.03 2.5 7.03 2.96 0.875 2.96  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.5585 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.585 3.19 17.945 3.19 17.945 1.475 10.27 1.475 10.27 1.14 10.61 1.14 10.61 1.245 12.51 1.245 12.51 1.14 15.09 1.14 15.09 1.245 16.99 1.245 16.99 1.14 18.175 1.14 18.175 3.45 18.33 3.45 18.33 3.83 16.205 3.83 16.205 4.36 15.975 4.36 15.975 3.42 11.625 3.42 11.625 4.36 11.395 4.36 11.395 3.42 7.095 3.42 7.095 4.36 6.865 4.36 6.865 3.42 2.815 3.42 2.815 4.36 2.585 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 4.675 4.59 4.675 3.65 4.905 3.65 4.905 4.59 9.105 4.59 9.105 3.65 9.335 3.65 9.335 4.59 13.635 4.59 13.635 3.65 13.865 3.65 13.865 4.59 18.065 4.59 18.065 4.06 18.295 4.06 18.295 4.59 18.635 4.59 19.04 4.59 19.04 5.49 18.635 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 8.315 0.45 8.315 1.07 8.085 1.07 8.085 0.45 6.075 0.45 6.075 1.07 5.845 1.07 5.845 0.45 3.835 0.45 3.835 1.07 3.605 1.07 3.605 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.73 0.475 0.73 0.475 1.31 2.485 1.31 2.485 0.73 2.715 0.73 2.715 1.31 4.725 1.31 4.725 0.73 4.955 0.73 4.955 1.31 6.965 1.31 6.965 0.73 7.195 0.73 7.195 1.31 9.205 1.31 9.205 0.68 18.635 0.68 18.635 1.54 18.405 1.54 18.405 0.91 16.21 0.91 16.21 1.015 15.87 1.015 15.87 0.91 11.73 0.91 11.73 1.015 11.39 1.015 11.39 0.91 9.435 0.91 9.435 1.54 0.245 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.135 1.77 2.135 2.555 1.83 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 1.77 3.26 1.77 3.26 2.5 2.92 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.99 1.77 4.33 1.77 4.33 2.5 3.99 2.5  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.77 0.97 1.77 0.97 2.5 0.63 2.5  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.5256 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.465 3.45 2.42 3.45 2.42 1.14 2.77 1.14 2.77 1.31 3.835 1.31 4.725 1.31 4.725 0.73 4.955 0.73 4.955 1.54 3.835 1.54 2.65 1.54 2.65 3.83 1.695 3.83 1.695 4.36 1.465 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 3.835 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 5.6 4.59 5.6 5.49 3.835 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 0.475 0.45 0.475 1.54 0.245 1.54 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.68 3.835 0.68 3.835 1.07 3.605 1.07 3.605 0.91 1.595 0.91 1.595 1.54 1.365 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 2.27 5.5 2.27 5.5 2.71 4.63 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 3.77 1.77 3.77 1.81 6.275 1.81 6.275 2.215 7.685 2.215 7.685 2.555 6.045 2.555 6.045 2.04 4.38 2.04 4.38 2.5 4.04 2.5 4.04 2.15 3.51 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.055 2.215 3.285 2.215 3.285 2.94 7.99 2.94 7.99 2.215 8.755 2.215 8.755 2.71 8.22 2.71 8.22 3.17 3.055 3.17  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.675 2.215 0.97 2.215 0.97 2.71 0.675 2.71  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.13145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.4 8.985 3.4 8.985 1.935 6.505 1.935 6.505 1.58 3.935 1.58 3.935 1.54 3.605 1.54 3.605 1.14 4.065 1.14 4.065 1.35 5.845 1.35 5.845 1.14 6.735 1.14 6.735 1.705 7.43 1.705 7.43 1.14 8.315 1.14 8.315 1.705 9.215 1.705 9.215 3.63 6.025 3.63 6.025 4.36 5.795 4.36 5.795 3.63 1.595 3.63 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.86 0.525 3.86 0.525 4.59 2.385 4.59 2.385 3.86 2.615 3.86 2.615 4.59 9.105 4.59 9.105 3.86 9.335 3.86 9.335 4.59 9.67 4.59 10.08 4.59 10.08 5.49 9.67 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 1.595 0.45 1.595 1.525 1.365 1.525 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.755 2.485 1.755 2.485 0.68 9.67 0.68 9.67 1.655 9.44 1.655 9.44 0.91 7.195 0.91 7.195 1.185 6.965 1.185 6.965 0.91 4.955 0.91 4.955 1.12 4.725 1.12 4.725 0.91 2.715 0.91 2.715 1.985 0.245 1.985  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.59 2.27 7.99 2.27 7.99 1.77 10.39 1.77 10.39 2.27 11.1 2.27 11.1 2.5 10.16 2.5 10.16 2 8.25 2 8.25 2.5 7.59 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.355 2.215 5.585 2.215 5.585 2.73 9.59 2.73 9.59 2.27 9.93 2.27 9.93 2.73 13.005 2.73 13.005 2.215 13.235 2.215 13.235 2.96 5.355 2.96  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.77 1.53 1.77 1.53 2.27 3.89 2.27 3.89 2.5 1.27 2.5  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.27 2.27 17.85 2.27 17.85 2.71 15.27 2.71  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.50965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.96 3.605 11.395 3.605 11.395 3.19 13.465 3.19 13.465 1.985 10.62 1.985 10.62 1.54 7.825 1.54 7.825 1.605 1.695 1.605 1.695 1.54 1.365 1.54 1.365 1.14 1.86 1.14 1.86 1.375 3.55 1.375 3.55 1.14 3.89 1.14 3.89 1.375 5.19 1.375 5.19 1.14 6.13 1.14 6.13 1.375 7.66 1.375 7.66 1.14 8.37 1.14 8.37 1.31 10.27 1.31 10.27 1.14 10.85 1.14 10.85 1.755 12.565 1.755 12.565 1.14 12.795 1.14 12.795 1.755 13.695 1.755 13.695 3.09 17.745 3.09 17.745 4.36 17.515 4.36 17.515 3.32 15.555 3.32 15.555 4.36 15.325 4.36 15.325 3.42 11.625 3.42 11.625 3.89 6.96 3.89  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.55 1.595 3.55 1.595 4.59 3.555 4.59 3.555 3.55 3.785 3.55 3.785 4.59 13.87 4.59 14.305 4.59 14.305 3.875 14.535 3.875 14.535 4.59 16.495 4.59 16.495 3.55 16.725 3.55 16.725 4.59 18.635 4.59 18.635 3.55 18.865 3.55 18.865 4.59 18.915 4.59 19.6 4.59 19.6 5.49 18.915 5.49 13.87 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.6 -0.45 19.6 0.45 17.795 0.45 17.795 1.58 17.565 1.58 17.565 0.45 15.555 0.45 15.555 1.58 15.325 1.58 15.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 3.09 5.165 3.09 5.165 4.12 13.87 4.12 13.87 4.35 4.935 4.35 4.935 3.32 2.715 3.32 2.715 4.36 2.485 4.36 2.485 3.32 0.575 3.32 0.575 4.36 0.345 4.36  ;
        POLYGON 0.245 0.68 14.155 0.68 14.155 1.81 16.445 1.81 16.445 0.805 16.675 0.805 16.675 1.81 18.685 1.81 18.685 0.805 18.915 0.805 18.915 2.04 13.925 2.04 13.925 0.91 11.675 0.91 11.675 1.525 11.445 1.525 11.445 0.91 9.49 0.91 9.49 1.08 9.15 1.08 9.15 0.91 7.195 0.91 7.195 1.145 6.965 1.145 6.965 0.91 4.955 0.91 4.955 1.145 4.725 1.145 4.725 0.91 2.715 0.91 2.715 1.145 2.485 1.145 2.485 0.91 0.475 0.91 0.475 1.615 0.245 1.615  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.72 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.555 4.07 2.555  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 1.77 5.45 1.77 5.45 2.555 5.19 2.555  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.655 2.785 4.63 2.785 4.63 1.14 4.955 1.14 4.955 3.015 3.885 3.015 3.885 4.36 3.655 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 5.745 4.59 5.745 3.55 5.975 3.55 5.975 4.59 6.075 4.59 6.72 4.59 6.72 5.49 6.075 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.72 -0.45 6.72 0.45 2.715 0.45 2.715 1.58 2.485 1.58 2.485 0.45 0.475 0.45 0.475 1.58 0.245 1.58 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.77 1.595 0.77 1.595 1.81 3.605 1.81 3.605 0.68 6.075 0.68 6.075 1.58 5.845 1.58 5.845 0.91 3.835 0.91 3.835 2.04 1.365 2.04  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 2.27 2.46 2.27 2.46 1.81 4.63 1.81 4.63 1.77 4.89 1.77 4.89 2.27 5.45 2.27 5.45 2.5 4.63 2.5 4.63 2.04 2.69 2.04 2.69 2.5 1.94 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.94 5.68 2.94 5.68 2.27 6.57 2.27 6.57 2.5 5.91 2.5 5.91 3.17 0.71 3.17  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.515 2.215 8.81 2.215 8.81 2.71 8.515 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 2.215 7.735 2.215 7.735 2.94 10.765 2.94 10.765 2.215 10.995 2.215 10.995 3.17 7.43 3.17  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.655 3.415 11.225 3.415 11.225 1.985 7.99 1.985 7.99 1.14 8.315 1.14 8.315 1.755 10.325 1.755 10.325 1.14 10.555 1.14 10.555 1.755 11.455 1.755 11.455 3.645 9.385 3.645 9.385 4.34 9.155 4.34 9.155 3.645 3.885 3.645 3.885 4.355 3.655 4.355  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.875 0.575 3.875 0.575 4.59 6.865 4.59 6.865 3.875 7.095 3.875 7.095 4.59 11.345 4.59 11.345 3.875 11.575 3.875 11.575 4.59 11.915 4.59 12.32 4.59 12.32 5.49 11.915 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 6.075 0.45 6.075 1.095 5.845 1.095 5.845 0.45 3.835 0.45 3.835 1.095 3.605 1.095 3.605 0.45 1.595 0.45 1.595 1.095 1.365 1.095 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.755 0.475 0.755 0.475 1.335 2.485 1.335 2.485 0.755 2.715 0.755 2.715 1.335 4.37 1.335 4.37 1.31 4.725 1.31 4.725 0.73 5.16 0.73 5.16 1.335 6.965 1.335 6.965 0.68 11.915 0.68 11.915 1.565 11.685 1.565 11.685 0.91 9.435 0.91 9.435 1.525 9.205 1.525 9.205 0.91 7.195 0.91 7.195 1.565 5.055 1.565 5.055 1.54 4.475 1.54 4.475 1.565 0.245 1.565  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.67 2.27 13.055 2.27 13.055 2.71 9.67 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.08 2.215 1.31 2.215 1.31 2.785 4.245 2.785 4.245 2.27 7.13 2.27 7.13 2.785 8.78 2.785 8.78 2.215 9.01 2.215 9.01 3.015 6.87 3.015 6.87 2.5 4.475 2.5 4.475 3.015 1.08 3.015  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.37 1.81 7.43 1.81 7.43 1.77 7.69 1.77 7.69 2.555 7.43 2.555 7.43 2.04 3.6 2.04 3.6 2.555 3.37 2.555  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.275 1.81 20.31 1.81 20.31 1.77 20.57 1.77 20.57 2.27 20.785 2.27 20.785 2.5 20.31 2.5 20.31 2.04 17.615 2.04 17.615 2.5 17.275 2.5  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.035 2.27 15.535 2.27 15.535 2.73 17.845 2.73 17.845 2.27 18.86 2.27 18.86 2.73 22.36 2.73 22.36 2.215 22.59 2.215 22.59 2.96 18.89 2.96 18.89 3.27 18.63 3.27 18.63 2.5 18.075 2.5 18.075 2.96 15.305 2.96 15.305 2.5 15.035 2.5  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.467 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.53 3.09 15.115 3.09 15.115 3.19 16.93 3.19 16.93 3.45 17.21 3.45 17.21 3.77 21.08 3.77 21.08 3.19 22.82 3.19 22.82 1.565 20.675 1.565 20.675 1.54 20.07 1.54 20.07 1.57 15.53 1.57 15.53 1.14 15.76 1.14 15.76 1.34 17.77 1.34 17.77 1.14 18 1.14 18 1.34 19.955 1.34 19.955 1.14 20.78 1.14 20.78 1.335 22.25 1.335 22.25 1.14 23.05 1.14 23.05 3.42 21.31 3.42 21.31 4 16.7 4 16.7 3.42 14.925 3.42 14.925 3.32 12.8 3.32 12.8 3.9 12.57 3.9 12.57 3.32 10.76 3.32 10.76 3.9 10.53 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.59 4.59 2.59 3.705 2.82 3.705 2.82 4.59 7.07 4.59 7.07 3.705 7.3 3.705 7.3 4.59 14.02 4.59 14.51 4.59 14.51 3.56 14.74 3.56 14.74 4.59 18.84 4.59 18.84 4.345 19.07 4.345 19.07 4.59 23.28 4.59 23.28 3.09 23.51 3.09 23.51 4.59 23.6 4.59 24.08 4.59 24.08 5.49 23.6 5.49 14.02 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 24.08 -0.45 24.08 0.45 13 0.45 13 1.11 12.77 1.11 12.77 0.45 10.76 0.45 10.76 1.11 10.53 1.11 10.53 0.45 8.52 0.45 8.52 1.11 8.29 1.11 8.29 0.45 6.28 0.45 6.28 1.11 6.05 1.11 6.05 0.45 4.04 0.45 4.04 1.11 3.81 1.11 3.81 0.45 1.8 0.45 1.8 1.11 1.57 1.11 1.57 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.5 3.09 0.73 3.09 0.73 3.245 4.88 3.245 4.88 3.09 5.11 3.09 5.11 3.245 7.76 3.245 7.76 4.13 11.55 4.13 11.55 3.55 11.78 3.55 11.78 4.13 13.79 4.13 13.79 3.55 14.02 3.55 14.02 4.36 7.53 4.36 7.53 3.475 5.11 3.475 5.11 3.9 4.88 3.9 4.88 3.475 0.73 3.475 0.73 3.9 0.5 3.9  ;
        POLYGON 0.45 0.77 0.68 0.77 0.68 1.35 2.69 1.35 2.69 0.77 2.92 0.77 2.92 1.35 4.93 1.35 4.93 0.77 5.16 0.77 5.16 1.35 7.17 1.35 7.17 0.73 7.4 0.73 7.4 1.31 7.95 1.31 7.95 1.35 9.41 1.35 9.41 0.77 9.64 0.77 9.64 1.35 11.65 1.35 11.65 0.77 11.88 0.77 11.88 1.35 13.89 1.35 13.89 0.68 23.6 0.68 23.6 1.58 23.37 1.58 23.37 0.91 21.36 0.91 21.36 1.105 21.13 1.105 21.13 0.91 19.12 0.91 19.12 1.11 18.89 1.11 18.89 0.91 16.88 0.91 16.88 1.11 16.65 1.11 16.65 0.91 14.12 0.91 14.12 1.58 7.82 1.58 7.82 1.54 7.3 1.54 7.3 1.58 0.45 1.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.555 4.07 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 2.215 5.45 2.215 5.45 3.27 5.19 3.27  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.23 2.27 6.57 2.27 6.57 2.71 6.23 2.71  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.4018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.655 2.785 4.67 2.785 4.67 1.14 4.955 1.14 4.955 1.755 6.075 1.755 6.31 1.755 6.31 1.21 6.965 1.21 6.965 0.715 7.195 0.715 7.195 1.59 6.54 1.59 6.54 1.985 6.075 1.985 4.9 1.985 4.9 3.015 3.885 3.015 3.885 4.36 3.655 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 6.075 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 7.84 4.59 7.84 5.49 6.075 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 2.715 0.45 2.715 1.525 2.485 1.525 2.485 0.45 0.475 0.45 0.475 1.525 0.245 1.525 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.715 1.595 0.715 1.595 1.755 2.945 1.755 2.945 0.68 6.075 0.68 6.075 1.525 5.845 1.525 5.845 0.91 3.835 0.91 3.835 1.525 3.605 1.525 3.605 0.91 3.175 0.91 3.175 1.985 1.365 1.985  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.59 2.28 9.93 2.28 9.93 2.71 9.59 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.55 1.77 8.81 1.77 8.81 1.82 10.39 1.82 10.39 2.27 12.22 2.27 12.22 2.5 10.16 2.5 10.16 2.05 8.89 2.05 8.89 2.5 8.55 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 2.215 7.735 2.215 7.735 2.94 13.005 2.94 13.005 2.215 13.235 2.215 13.235 3.17 7.43 3.17  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.99 2.27 2.39 2.27 2.39 1.77 3.72 1.77 3.72 2.27 5.5 2.27 5.5 2.5 3.49 2.5 3.49 2 2.65 2 2.65 2.5 1.99 2.5  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.94 5.73 2.94 5.73 2.27 6.62 2.27 6.62 2.5 5.96 2.5 5.96 3.17 0.71 3.17  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.3284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.655 3.4 13.465 3.4 13.465 1.59 10.23 1.59 10.23 1.48 8.03 1.48 8.03 1.25 10.23 1.25 10.23 1.14 10.555 1.14 10.555 1.25 13.695 1.25 13.695 3.63 10.505 3.63 10.505 4.36 10.275 4.36 10.275 3.63 3.885 3.63 3.885 4.36 3.655 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.86 0.575 3.86 0.575 4.59 6.915 4.59 6.915 3.86 7.145 3.86 7.145 4.59 13.585 4.59 13.585 3.86 13.815 3.86 13.815 4.59 13.915 4.59 14.56 4.59 14.56 5.49 13.915 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 6.075 0.45 6.075 1.565 5.845 1.565 5.845 0.45 3.835 0.45 3.835 1 3.605 1 3.605 0.45 1.595 0.45 1.595 1.455 1.365 1.455 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.685 1.93 1.685 1.93 0.73 2.715 0.73 2.715 1.31 4.725 1.31 4.725 0.73 4.955 0.73 4.955 1.795 6.965 1.795 6.965 0.68 13.915 0.68 13.915 1.02 11.445 1.02 11.445 0.91 9.435 0.91 9.435 1.02 7.195 1.02 7.195 2.025 4.725 2.025 4.725 1.54 2.16 1.54 2.16 1.915 0.245 1.915  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 28.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.325 2.19 17.85 2.19 17.85 2.71 15.325 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.12 2.27 19.46 2.27 19.46 2.495 21.99 2.495 21.99 2.27 22.82 2.27 22.82 2.495 26.965 2.495 26.965 2.215 27.195 2.215 27.195 2.725 19.12 2.725  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.69 1.81 25.06 1.81 25.06 2.265 24.72 2.265 24.72 2.04 20.58 2.04 20.58 2.265 19.69 2.265  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.325 2.19 12.795 2.19 12.795 2.71 10.325 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.82 2.19 1.16 2.19 1.16 2.65 4.04 2.65 4.04 2.27 4.38 2.27 4.38 2.65 6.8 2.65 6.8 2.27 8.86 2.27 8.86 2.5 7.03 2.5 7.03 2.88 0.82 2.88  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 4.84 1.77 4.84 2.19 6.57 2.19 6.57 2.42 4.61 2.42 4.61 2 2.17 2 2.17 2.42 1.83 2.42  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.3823 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.325 2.955 27.425 2.955 27.425 1.53 15.27 1.53 15.27 1.3 17.51 1.3 17.51 1.14 17.85 1.14 17.85 1.3 19.75 1.3 19.75 1.14 20.09 1.14 20.09 1.3 21.99 1.3 21.99 1.14 22.33 1.14 22.33 1.3 24.23 1.3 24.23 1.14 24.57 1.14 24.57 1.3 27.655 1.3 27.655 3.185 17.745 3.185 17.745 3.46 17.515 3.46 17.515 3.185 15.555 3.185 15.555 3.46 15.325 3.46 15.325 3.185 13.85 3.185 13.85 3.83 12.565 3.83 12.565 3.185 10.555 3.185 10.555 3.83 10.325 3.83  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.58 2.615 3.58 2.615 4.59 6.865 4.59 6.865 3.58 7.095 3.58 7.095 4.59 13.87 4.59 20.875 4.59 20.875 4.15 21.105 4.15 21.105 4.59 25.355 4.59 25.355 3.875 25.585 3.875 25.585 4.59 27.775 4.59 27.875 4.59 28.56 4.59 28.56 5.49 27.875 5.49 27.775 5.49 13.87 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 28.56 -0.45 28.56 0.45 12.795 0.45 12.795 1.07 12.565 1.07 12.565 0.45 10.555 0.45 10.555 1.07 10.325 1.07 10.325 0.45 8.315 0.45 8.315 1.07 8.085 1.07 8.085 0.45 6.075 0.45 6.075 1.07 5.845 1.07 5.845 0.45 3.835 0.45 3.835 1.07 3.605 1.07 3.605 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 3.12 7.555 3.12 7.555 4.06 11.345 4.06 11.345 3.48 11.575 3.48 11.575 4.06 13.87 4.06 13.87 4.29 7.325 4.29 7.325 3.35 4.905 3.35 4.905 3.93 4.675 3.93 4.675 3.35 0.525 3.35 0.525 3.93 0.295 3.93  ;
        POLYGON 14.305 3.48 14.535 3.48 14.535 3.69 16.445 3.69 16.445 3.48 16.675 3.48 16.675 3.69 23.115 3.69 23.115 3.415 27.775 3.415 27.775 4.225 27.545 4.225 27.545 3.645 23.345 3.645 23.345 3.92 14.305 3.92  ;
        POLYGON 0.245 0.73 0.475 0.73 0.475 1.31 2.485 1.31 2.485 0.73 2.715 0.73 2.715 1.31 4.725 1.31 4.725 0.73 4.955 0.73 4.955 1.31 6.965 1.31 6.965 0.73 7.195 0.73 7.195 1.31 9.205 1.31 9.205 0.73 9.435 0.73 9.435 1.31 11.445 1.31 11.445 0.73 11.675 0.73 11.675 1.31 14.2 1.31 14.2 0.68 27.875 0.68 27.875 1.07 25.405 1.07 25.405 0.91 23.45 0.91 23.45 1.015 23.11 1.015 23.11 0.91 21.21 0.91 21.21 1.015 20.87 1.015 20.87 0.91 18.97 0.91 18.97 1.015 18.63 1.015 18.63 0.91 16.675 0.91 16.675 1.07 14.43 1.07 14.43 1.54 0.245 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.27 2.17 2.27 2.17 2.71 1.83 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.27 3.29 2.27 3.29 2.71 2.95 2.71  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.99 2.27 4.33 2.27 4.33 2.71 3.99 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.4988 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.14 1.595 1.14 1.595 3.09 2.715 3.09 4.835 3.09 4.835 4.36 4.605 4.36 4.605 3.32 2.715 3.32 2.615 3.32 2.615 4.36 2.385 4.36 2.385 3.32 1.27 3.32  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 2.715 4.59 3.585 4.59 3.585 3.55 3.815 3.55 3.815 4.59 5.6 4.59 5.6 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.835 0.45 4.835 1.655 4.605 1.655 4.605 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 2.715 0.68 2.715 1.655 2.485 1.655 2.485 0.91 0.475 0.91 0.475 1.655 0.245 1.655  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.795 2.215 2.09 2.215 2.09 2.71 1.795 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 2.27 1.54 2.27 1.54 2.94 2.39 2.94 2.39 2.27 4.33 2.27 4.33 2.71 2.62 2.71 2.62 3.17 1.2 3.17  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.33 2.27 5.67 2.27 5.67 2.94 6.87 2.94 6.87 2.215 8.535 2.215 8.535 3.17 5.33 3.17  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.23 2.27 6.57 2.27 6.57 2.71 6.23 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.0258 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 3.375 1.095 3.375 1.095 4.07 2.435 4.07 2.435 3.4 8.095 3.4 8.095 4.36 7.865 4.36 7.865 3.63 6.055 3.63 6.055 4.36 5.825 4.36 5.825 3.63 2.665 3.63 2.665 4.36 0.865 4.36 0.865 3.58 0.74 3.58 0.74 1.14 1.595 1.14 1.595 1.34 3.89 1.34 3.89 1.57 0.97 1.57  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.86 0.575 3.86 0.575 4.59 4.625 4.59 4.625 3.86 4.855 3.86 4.855 4.59 6.845 4.59 6.845 3.86 7.075 3.86 7.075 4.59 8.885 4.59 8.885 3.86 9.115 3.86 9.115 4.59 9.52 4.59 9.52 5.49 9.115 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 7.075 0.45 7.075 1.525 6.845 1.525 6.845 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 4.955 0.68 4.955 1.755 8.885 1.755 8.885 0.77 9.115 0.77 9.115 1.985 4.725 1.985 4.725 1.11 2.485 1.11 2.485 0.91 0.475 0.91 0.475 1.58 0.245 1.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.06 2.39 3.51 2.39 3.51 1.77 3.77 1.77 3.77 1.87 4.79 1.87 4.79 2.39 6.62 2.39 6.62 2.62 4.56 2.62 4.56 2.1 3.77 2.1 3.77 2.62 3.06 2.62  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.39 1.21 2.39 1.21 2.85 4.07 2.85 4.07 2.33 4.33 2.33 4.33 2.85 6.85 2.85 6.85 2.39 8.81 2.39 8.81 2.62 7.08 2.62 7.08 3.08 0.87 3.08  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.67 2.33 9.955 2.33 9.955 2.85 12.875 2.85 12.875 2.335 13.105 2.335 13.105 2.85 15.24 2.85 15.24 2.39 17.15 2.39 17.15 2.62 15.47 2.62 15.47 3.08 9.67 3.08  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.85 2.39 12.27 2.39 12.27 2 12.33 2 12.33 1.77 13.565 1.77 13.565 2.39 15.01 2.39 15.01 2.62 13.335 2.62 13.335 2 12.73 2 12.73 2.155 12.5 2.155 12.5 2.62 11.85 2.62  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.9601 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.64 3.31 16.655 3.31 16.655 4.36 16.425 4.36 16.425 3.54 14.615 3.54 14.615 4.345 14.385 4.345 14.385 3.54 12.575 3.54 12.575 4.36 12.345 4.36 12.345 3.83 11.91 3.83 11.91 3.54 10.535 3.54 10.535 4.12 10.305 4.12 10.305 3.54 7.145 3.54 7.145 4.36 6.915 4.36 6.915 3.54 2.715 3.54 2.715 4.36 2.485 4.36 2.485 3.54 0.41 3.54 0.41 1.72 1.365 1.72 1.365 1.14 1.595 1.14 1.595 1.72 3.05 1.72 3.05 1.14 4.12 1.14 4.12 1.35 5.845 1.35 5.845 1.14 6.21 1.14 6.21 1.6 8.085 1.6 8.085 1.14 8.315 1.14 8.315 1.83 5.98 1.83 5.98 1.58 3.99 1.58 3.99 1.54 3.28 1.54 3.28 1.95 0.64 1.95  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.77 0.575 3.77 0.575 4.59 4.675 4.59 4.675 3.77 4.905 3.77 4.905 4.59 9.105 4.59 9.105 3.77 9.335 3.77 9.335 4.59 11.325 4.59 11.325 3.77 11.555 3.77 11.555 4.59 13.365 4.59 13.365 3.77 13.595 3.77 13.595 4.59 15.405 4.59 15.405 3.77 15.635 3.77 15.635 4.59 17.445 4.59 17.445 3.77 17.675 3.77 17.675 4.59 17.92 4.59 17.92 5.49 17.675 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 15.635 0.45 15.635 1.49 15.405 1.49 15.405 0.45 11.555 0.45 11.555 1.265 11.325 1.265 11.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 9.435 0.68 9.435 1.495 11.87 1.495 11.87 1.31 13.365 1.31 13.365 0.68 13.595 0.68 13.595 1.31 14.025 1.31 14.025 1.72 17.445 1.72 17.445 0.68 17.675 0.68 17.675 1.95 13.795 1.95 13.795 1.54 12.1 1.54 12.1 1.725 9.205 1.725 9.205 0.91 7.25 0.91 7.25 0.965 6.91 0.965 6.91 0.91 5.01 0.91 5.01 0.965 4.67 0.965 4.67 0.91 2.77 0.91 2.77 0.965 2.43 0.965 2.43 0.91 0.475 0.91 0.475 1.49 0.245 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.72 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 1.77 5.455 1.77 5.455 2.555 5.19 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 2.215 4.435 2.215 4.435 2.71 4.07 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.15 2.09 2.15 2.09 2.71 1.83 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.015 1.77 1.015 2.555 0.71 2.555  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.27 3.29 2.27 3.29 2.71 2.95 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.6616 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.895 3.09 6.035 3.09 6.035 4.36 5.805 4.36 5.805 3.32 2.795 3.32 2.795 4.36 2.715 4.36 2.565 4.36 2.565 3.09 2.715 3.09 4.665 3.09 4.665 1.59 4.63 1.59 4.63 1.14 5.015 1.14 5.015 1.48 4.895 1.48  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 2.715 4.59 3.585 4.59 3.585 3.55 3.815 3.55 3.815 4.59 6.135 4.59 6.72 4.59 6.72 5.49 6.135 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.72 -0.45 6.72 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.73 0.475 0.73 0.475 1.31 2.485 1.31 2.485 0.73 2.715 0.73 2.715 1.54 0.245 1.54  ;
        POLYGON 3.665 0.68 6.135 0.68 6.135 1.54 5.905 1.54 5.905 0.91 3.895 0.91 3.895 1.54 3.665 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.53 2.215 7.76 2.215 7.76 2.89 9.075 2.89 9.075 2.27 11.14 2.27 11.14 2.5 9.305 2.5 9.305 3.27 7.53 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.99 1.77 8.25 1.77 8.25 2.215 8.845 2.215 8.845 2.555 7.99 2.555  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.15 3.21 2.15 3.21 2.71 2.95 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 1.83 2.165 1.83 2.165 2.325 2.5 2.325 2.5 2.94 4.575 2.94 4.575 2.215 5.425 2.215 5.425 2.555 4.805 2.555 4.805 3.17 2.27 3.17 2.27 2.555 1.21 2.555  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 3.35 2.125 3.35 2.125 3.4 5.035 3.4 5.035 2.785 6.16 2.785 6.395 2.785 6.395 2.215 6.625 2.215 6.625 3.015 6.16 3.015 5.265 3.015 5.265 3.63 1.98 3.63 1.98 3.58 0.71 3.58  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.2165 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.295 3.81 1.835 3.81 1.835 3.86 5.495 3.86 5.495 3.55 6.16 3.55 10.79 3.55 10.79 2.89 11.435 2.89 11.435 1.985 8.48 1.985 8.48 1.54 8.12 1.54 8.12 1.31 8.71 1.31 8.71 1.755 10.415 1.755 10.415 1.14 10.645 1.14 10.645 1.755 11.665 1.755 11.665 3.78 7.205 3.78 7.205 4.36 6.975 4.36 6.975 3.78 6.16 3.78 5.725 3.78 5.725 4.09 3.765 4.09 3.765 4.36 3.535 4.36 3.535 4.09 1.69 4.09 1.69 4.04 0.525 4.04 0.525 4.36 0.295 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 4.27 1.545 4.27 1.545 4.59 5.955 4.59 5.955 4.02 6.16 4.02 6.185 4.02 6.185 4.59 9.245 4.59 9.245 4.02 9.475 4.02 9.475 4.59 11.765 4.59 12.32 4.59 12.32 5.49 11.765 5.49 6.16 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 5.04 0.45 5.04 0.64 4.7 0.64 4.7 0.45 2.8 0.45 2.8 0.64 2.46 0.64 2.46 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.34 1.33 6.16 1.33 6.16 1.56 1.34 1.56  ;
        POLYGON 0.245 0.715 0.475 0.715 0.475 0.87 7.055 0.87 7.055 0.68 11.765 0.68 11.765 1.525 11.535 1.525 11.535 0.91 9.525 0.91 9.525 1.525 9.295 1.525 9.295 0.91 7.285 0.91 7.285 1.19 7.055 1.19 7.055 1.1 0.475 1.1 0.475 1.525 0.245 1.525  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.03 2.27 15.37 2.27 15.37 3.04 19.14 3.04 19.14 2.215 19.37 2.215 19.37 2.89 20.96 2.89 20.96 2.27 22.97 2.27 22.97 2.5 21.19 2.5 21.19 3.27 15.03 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.27 2.27 17.51 2.27 17.51 1.755 19.83 1.755 19.83 2.27 20.73 2.27 20.73 2.5 19.6 2.5 19.6 1.985 17.77 1.985 17.77 2.5 17.27 2.5  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.27 1.21 2.27 1.21 2.73 4.07 2.73 4.07 2.27 4.41 2.27 4.41 2.73 6.85 2.73 6.85 2.27 8.86 2.27 8.86 2.5 7.08 2.5 7.08 2.96 0.87 2.96  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.06 2.27 3.4 2.27 3.4 2.02 3.46 2.02 3.46 1.77 4.87 1.77 4.87 2.27 6.62 2.27 6.62 2.5 4.64 2.5 4.64 2.04 3.86 2.04 3.86 2.175 3.63 2.175 3.63 2.5 3.06 2.5  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.99 2.27 13.515 2.27 13.57 2.27 13.57 2.71 13.515 2.71 10.99 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.615 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.345 3.19 4.905 3.19 4.905 3.5 13.515 3.5 23.2 3.5 23.2 1.97 20.06 1.97 20.06 1.52 15.525 1.52 15.525 1.14 15.755 1.14 15.755 1.29 17.71 1.29 17.71 1.14 18.05 1.14 18.05 1.29 20.005 1.29 20.005 1.14 20.29 1.14 20.29 1.74 22.245 1.74 22.245 1.14 22.475 1.14 22.475 1.74 23.495 1.74 23.495 4.36 23.265 4.36 23.265 3.73 19.065 3.73 19.065 4.36 18.57 4.36 18.57 3.73 14.535 3.73 14.535 4.36 14.305 4.36 14.305 3.73 13.515 3.73 12.395 3.73 12.395 4.36 12.165 4.36 12.165 3.73 9.385 3.73 9.385 4.36 9.155 4.36 9.155 3.73 4.905 3.73 4.905 4.36 4.675 4.36 4.675 3.42 0.575 3.42 0.575 4.36 0.345 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.65 2.665 3.65 2.665 4.59 6.915 4.59 6.915 3.96 7.145 3.96 7.145 4.59 10.945 4.59 10.945 3.96 11.175 3.96 11.175 4.59 13.185 4.59 13.185 3.96 13.415 3.96 13.415 4.59 13.515 4.59 16.595 4.59 16.595 3.96 16.825 3.96 16.825 4.59 21.075 4.59 21.075 3.96 21.305 3.96 21.305 4.59 23.595 4.59 24.08 4.59 24.08 5.49 23.595 5.49 13.515 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 24.08 -0.45 24.08 0.45 9.435 0.45 9.435 1.04 9.205 1.04 9.205 0.45 7.195 0.45 7.195 1.04 6.965 1.04 6.965 0.45 4.955 0.45 4.955 1.04 4.725 1.04 4.725 0.45 2.715 0.45 2.715 1.51 2.485 1.51 2.485 0.45 0.475 0.45 0.475 1.51 0.245 1.51 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.7 1.595 0.7 1.595 1.74 2.945 1.74 2.945 1.28 3.605 1.28 3.605 0.7 3.835 0.7 3.835 1.28 5.845 1.28 5.845 0.7 6.075 0.7 6.075 1.28 8.085 1.28 8.085 0.7 8.315 0.7 8.315 1.28 10.99 1.28 10.99 1.14 11.33 1.14 11.33 1.28 13.285 1.28 13.285 1.14 13.515 1.14 13.515 1.51 3.175 1.51 3.175 1.97 1.365 1.97  ;
        POLYGON 9.925 0.68 23.595 0.68 23.595 1.51 23.365 1.51 23.365 0.91 21.355 0.91 21.355 1.51 21.125 1.51 21.125 0.91 19.17 0.91 19.17 0.985 18.83 0.985 18.83 0.91 16.93 0.91 16.93 0.985 16.59 0.985 16.59 0.91 14.69 0.91 14.69 0.985 14.35 0.985 14.35 0.91 12.45 0.91 12.45 0.985 12.11 0.985 12.11 0.91 10.155 0.91 10.155 1.04 9.925 1.04  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.4 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.87 2.27 7.29 2.27 7.29 2.71 6.87 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 2.27 6.18 2.27 6.18 2.71 5.75 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 3.98 1.77 3.98 2.5 3.51 2.5  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 2.27 5.05 2.27 5.05 2.71 4.63 2.71  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.15 2.09 2.15 2.09 2.71 1.83 2.71  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.9438 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.64 3.55 7.815 3.55 7.815 4.36 7.585 4.36 7.585 3.83 4.555 3.83 3.485 3.83 3.485 4.36 3.255 4.36 3.255 3.45 4.555 3.45 6.41 3.45 6.41 1.14 6.795 1.14 6.795 1.48 6.64 1.48  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 4.555 4.59 5.345 4.59 5.345 4.06 5.575 4.06 5.575 4.59 7.915 4.59 8.4 4.59 8.4 5.49 7.915 5.49 4.555 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.4 -0.45 8.4 0.45 2.715 0.45 2.715 1.205 2.485 1.205 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.68 1.595 0.68 1.595 1.435 3.1 1.435 3.1 1.31 4.325 1.31 4.325 1.14 4.555 1.14 4.555 1.54 3.305 1.54 3.305 1.665 1.365 1.665  ;
        POLYGON 3.15 0.68 7.915 0.68 7.915 1.49 7.685 1.49 7.685 0.91 5.675 0.91 5.675 1.49 5.445 1.49 5.445 0.91 3.49 0.91 3.49 0.965 3.15 0.965  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.12 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.605 2.215 10.835 2.215 10.835 2.94 12.27 2.94 12.27 2.215 14.005 2.215 14.005 2.71 12.5 2.71 12.5 3.17 10.605 3.17  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.35 2.215 11.715 2.215 11.715 2.71 11.35 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 2.215 6.165 2.215 6.165 3.04 9.035 3.04 9.295 3.04 9.295 2.215 9.525 2.215 9.525 3.27 9.035 3.27 5.19 3.27  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.87 2.215 7.285 2.215 7.285 2.71 6.87 2.71  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.925 2.215 1.155 2.215 1.155 2.785 4.07 2.785 4.07 1.77 4.33 1.77 4.33 3.015 0.925 3.015  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.57 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.345 3.32 4.9 3.32 4.9 3.5 8.87 3.5 8.87 4.13 9.035 4.13 9.875 4.13 9.875 3.4 14.355 3.4 14.355 1.95 11.045 1.95 11.045 1.14 11.275 1.14 11.275 1.72 13.285 1.72 13.285 1.14 13.515 1.14 13.515 1.72 14.585 1.72 14.585 4.36 14.355 4.36 14.355 3.63 10.105 3.63 10.105 4.36 9.035 4.36 8.49 4.36 8.49 3.73 4.905 3.73 4.905 4.36 4.675 4.36 4.675 3.55 0.575 3.55 0.575 4.36 0.345 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.78 2.665 3.78 2.665 4.59 7.635 4.59 7.635 3.96 7.865 3.96 7.865 4.59 9.035 4.59 12.115 4.59 12.115 3.86 12.345 3.86 12.345 4.59 14.635 4.59 15.12 4.59 15.12 5.49 14.635 5.49 9.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.12 -0.45 15.12 0.45 4.955 0.45 4.955 0.695 4.725 0.695 4.725 0.45 2.715 0.45 2.715 0.695 2.485 0.695 2.485 0.45 0.475 0.45 0.475 1.655 0.245 1.655 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.73 1.595 0.73 1.595 0.925 3.605 0.925 3.605 0.73 3.835 0.73 3.835 1.14 9.035 1.14 9.035 1.54 1.365 1.54  ;
        POLYGON 5.39 0.68 14.635 0.68 14.635 1.49 14.405 1.49 14.405 0.91 12.395 0.91 12.395 1.49 12.165 1.49 12.165 0.91 10.155 0.91 10.155 1.575 9.925 1.575 9.925 0.91 5.39 0.91  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 28.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.19 1.77 27.395 1.77 27.395 2.555 27.165 2.555 27.165 2 22.915 2 22.915 2.145 22.685 2.145 22.685 2 19.66 2 19.66 2.5 19.19 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.7 2.27 22.04 2.27 22.04 2.48 23.11 2.48 23.11 2.27 25.26 2.27 25.26 2.71 21.7 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.605 2.215 10.835 2.215 10.835 2.89 13.72 2.89 13.72 2.27 14.06 2.27 14.06 3.04 17.995 3.04 18.2 3.04 18.2 2.27 18.54 2.27 18.54 3.27 17.995 3.27 10.605 3.27  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.74 2.27 13.03 2.27 13.03 1.77 14.52 1.77 14.52 2.27 16.25 2.27 16.25 2.5 14.29 2.5 14.29 2 13.29 2 13.29 2.5 12.74 2.5  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.875 2.215 1.105 2.215 1.105 2.785 4.04 2.785 4.04 2.27 4.38 2.27 4.38 2.785 6.85 2.785 6.85 2.27 8.86 2.27 8.86 2.5 7.08 2.5 7.08 3.015 0.875 3.015  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.165 2.215 3.51 2.215 3.51 1.77 4.84 1.77 4.84 2.27 6.62 2.27 6.62 2.5 4.61 2.5 4.61 2 3.77 2 3.77 2.555 3.165 2.555  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.5296 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.295 3.245 9.38 3.245 9.38 3.5 17.995 3.5 18.835 3.5 18.835 3.09 27.745 3.09 27.745 1.515 20.005 1.515 20.005 1.14 20.235 1.14 20.235 1.285 22.19 1.285 22.19 1.14 22.53 1.14 22.53 1.285 24.43 1.285 24.43 1.14 24.77 1.14 24.77 1.285 26.67 1.285 26.67 1.14 27.01 1.14 27.01 1.285 27.975 1.285 27.975 4.36 27.745 4.36 27.745 3.32 23.495 3.32 23.495 4.36 23.265 4.36 23.265 3.32 19.065 3.32 19.065 4.36 18.835 4.36 18.835 3.73 17.995 3.73 14.585 3.73 14.585 4.36 12.97 4.36 12.97 3.73 9.385 3.73 9.385 4.36 9.155 4.36 9.155 3.55 4.905 3.55 4.905 4.36 4.675 4.36 4.675 3.475 0.525 3.475 0.525 4.36 0.295 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.705 2.665 3.705 2.665 4.59 6.915 4.59 6.915 3.78 7.145 3.78 7.145 4.59 12.115 4.59 12.115 3.96 12.345 3.96 12.345 4.59 16.595 4.59 16.595 3.96 16.825 3.96 16.825 4.59 17.995 4.59 21.075 4.59 21.075 3.55 21.305 3.55 21.305 4.59 25.555 4.59 25.555 3.55 25.785 3.55 25.785 4.59 28.075 4.59 28.56 4.59 28.56 5.49 28.075 5.49 17.995 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 28.56 -0.45 28.56 0.45 9.435 0.45 9.435 1.525 9.205 1.525 9.205 0.45 7.195 0.45 7.195 1.525 6.965 1.525 6.965 0.45 4.955 0.45 4.955 1.055 4.725 1.055 4.725 0.45 2.715 0.45 2.715 1.525 2.485 1.525 2.485 0.45 0.475 0.45 0.475 1.525 0.245 1.525 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.715 1.595 0.715 1.595 1.755 3.05 1.755 3.05 1.295 3.605 1.295 3.605 0.715 3.835 0.715 3.835 1.295 5.845 1.295 5.845 0.715 6.075 0.715 6.075 1.755 8.085 1.755 8.085 0.715 8.315 0.715 8.315 1.755 10.99 1.755 10.99 1.14 11.275 1.14 11.275 1.29 13.23 1.29 13.23 1.14 13.57 1.14 13.57 1.29 15.525 1.29 15.525 1.14 15.81 1.14 15.81 1.755 17.765 1.755 17.765 1.14 17.995 1.14 17.995 1.985 15.58 1.985 15.58 1.52 11.22 1.52 11.22 1.985 5.845 1.985 5.845 1.525 3.28 1.525 3.28 1.985 1.365 1.985  ;
        POLYGON 9.925 0.68 28.075 0.68 28.075 1.055 27.845 1.055 27.845 0.91 25.89 0.91 25.89 1 25.55 1 25.55 0.91 23.65 0.91 23.65 1 23.31 1 23.31 0.91 21.41 0.91 21.41 1 21.07 1 21.07 0.91 19.115 0.91 19.115 1.525 18.885 1.525 18.885 0.91 16.875 0.91 16.875 1.525 16.645 1.525 16.645 0.91 14.69 0.91 14.69 1 14.35 1 14.35 0.91 12.45 0.91 12.45 1 12.11 1 12.11 0.91 10.155 0.91 10.155 1.525 9.925 1.525  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.07 2.215 1.07 3.27 0.71 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.21 2.09 1.21 2.09 2.555 1.83 2.555  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.21 3.9 1.21 3.9 0.68 4.13 0.68 4.13 4.36 3.8 4.36 3.8 1.59 3.51 1.59  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.78 4.59 2.78 3.79 3.01 3.79 3.01 4.59 3.505 4.59 4.48 4.59 4.48 5.49 3.505 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 3.01 0.45 3.01 0.995 2.78 0.995 2.78 0.45 0.53 0.45 0.53 0.995 0.3 0.995 0.3 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 3.845 2.32 3.845 2.32 0.94 1.365 0.94 1.365 0.71 2.55 0.71 2.55 2.27 3.505 2.27 3.505 2.5 2.55 2.5 2.55 4.075 0.345 4.075  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.27 1.07 2.27 1.07 2.71 0.71 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.795 2.215 2.09 2.215 2.09 2.71 1.795 2.71  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 0.68 3.835 0.68 3.835 4.36 3.51 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.55 2.665 3.55 2.665 4.59 3.205 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 5.6 4.59 5.6 5.49 3.205 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 3.09 2.975 3.09 2.975 1.95 1.365 1.95 1.365 0.68 1.595 0.68 1.595 1.72 3.205 1.72 3.205 3.32 0.575 3.32 0.575 4.36 0.345 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.27 1.21 2.27 1.21 2.94 2.39 2.94 2.39 2.215 4.275 2.215 4.275 3.17 0.87 3.17  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5505 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.085 3.09 7.39 3.09 7.62 3.09 7.62 1.59 5.985 1.59 5.985 0.68 6.215 0.68 6.215 1.21 8.225 1.21 8.225 0.68 8.455 0.68 8.455 1.49 7.85 1.49 7.85 3.09 8.405 3.09 8.405 4.36 8.175 4.36 8.175 3.32 7.39 3.32 6.315 3.32 6.315 4.36 6.085 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 4.965 4.59 4.965 3.55 5.195 3.55 5.195 4.59 7.105 4.59 7.105 3.55 7.335 3.55 7.335 4.59 7.39 4.59 9.245 4.59 9.245 3.55 9.475 3.55 9.475 4.59 10.08 4.59 10.08 5.49 7.39 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 9.575 0.45 9.575 1.49 9.345 1.49 9.345 0.45 7.335 0.45 7.335 0.98 7.105 0.98 7.105 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.535 3.4 4.505 3.4 4.505 1.97 1.365 1.97 1.365 0.68 1.595 0.68 1.595 1.74 3.605 1.74 3.605 0.68 3.835 0.68 3.835 1.74 4.735 1.74 4.735 2.27 7.39 2.27 7.39 2.5 4.735 2.5 4.735 3.63 2.765 3.63 2.765 4.36 2.535 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.16 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7725 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 1.015 1.77 1.015 2.555 0.785 2.555 0.785 2.15 0.15 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7725 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7725 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.215 3.335 2.215 3.335 2.71 2.95 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.045 0.68 5.45 0.68 5.45 4.36 5.045 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 4.025 4.59 4.025 3.79 4.255 3.79 4.255 4.59 4.75 4.59 6.16 4.59 6.16 5.49 4.75 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.16 -0.45 6.16 0.45 4.015 0.45 4.015 0.86 3.785 0.86 3.785 0.45 1.595 0.45 1.595 0.86 1.365 0.86 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.29 3.845 3.565 3.845 3.565 1.32 0.245 1.32 0.245 0.68 0.475 0.68 0.475 1.09 2.485 1.09 2.485 0.68 2.715 0.68 2.715 1.09 3.795 1.09 3.795 2.27 4.75 2.27 4.75 2.5 3.795 2.5 3.795 4.075 0.29 4.075  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.72 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.27 1.07 2.27 1.07 2.71 0.71 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.795 2.215 2.09 2.215 2.09 2.71 1.795 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.915 2.215 3.21 2.215 3.21 2.71 2.915 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 2.89 4.905 2.89 4.905 0.68 5.135 0.68 5.135 4.36 4.63 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 3.555 4.59 3.555 3.55 3.785 3.55 3.785 4.59 4.505 4.59 5.925 4.59 5.925 3.55 6.155 3.55 6.155 4.59 6.72 4.59 6.72 5.49 4.505 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.72 -0.45 6.72 0.45 6.255 0.45 6.255 1.49 6.025 1.49 6.025 0.45 3.835 0.45 3.835 1.385 3.605 1.385 3.605 0.45 1.595 0.45 1.595 1.385 1.365 1.385 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 3.09 3.44 3.09 3.44 1.845 0.245 1.845 0.245 0.68 0.475 0.68 0.475 1.615 2.485 1.615 2.485 0.68 2.715 0.68 2.715 1.615 3.67 1.615 3.67 2.215 4.505 2.215 4.505 2.555 3.67 2.555 3.67 3.32 0.575 3.32 0.575 4.36 0.345 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.09 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.09 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 3.72 1.77 3.72 2.27 5.5 2.27 5.5 2.5 3.49 2.5 3.49 2 2.17 2 2.17 2.5 1.83 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.09 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.27 1.07 2.27 1.07 2.94 6.23 2.94 6.23 2.27 6.57 2.27 6.57 3.17 0.71 3.17  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.315 3.4 9.67 3.4 9.9 3.4 9.9 1.59 8.265 1.59 8.265 0.68 8.495 0.68 8.495 1.21 10.505 1.21 10.505 0.68 10.735 0.68 10.735 1.49 10.13 1.49 10.13 3.4 10.685 3.4 10.685 4.36 10.455 4.36 10.455 3.63 9.67 3.63 8.545 3.63 8.545 4.36 8.315 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.86 0.575 3.86 0.575 4.59 6.865 4.59 6.865 3.86 7.095 3.86 7.095 4.59 9.335 4.59 9.335 3.86 9.565 3.86 9.565 4.59 9.67 4.59 11.525 4.59 11.525 3.86 11.755 3.86 11.755 4.59 12.32 4.59 12.32 5.49 9.67 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 11.855 0.45 11.855 1.385 11.625 1.385 11.625 0.45 9.615 0.45 9.615 0.915 9.385 0.915 9.385 0.45 7.195 0.45 7.195 0.915 6.965 0.915 6.965 0.45 4.955 0.45 4.955 0.915 4.725 0.915 4.725 0.45 2.715 0.45 2.715 0.915 2.485 0.915 2.485 0.45 0.475 0.45 0.475 1.385 0.245 1.385 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 3.655 3.4 6.8 3.4 6.8 1.375 1.365 1.375 1.365 0.68 1.595 0.68 1.595 1.145 3.605 1.145 3.605 0.68 3.835 0.68 3.835 1.145 5.845 1.145 5.845 0.68 6.075 0.68 6.075 1.145 7.03 1.145 7.03 2.27 9.67 2.27 9.67 2.5 7.03 2.5 7.03 3.63 3.885 3.63 3.885 4.36 3.655 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6945 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 1.015 1.77 1.015 2.555 0.785 2.555 0.785 2.15 0.15 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6945 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.215 1.77 2.215 2.555 1.83 2.555  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6945 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.385 1.77 3.385 2.555 2.95 2.555  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6945 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.21 4.575 1.21 4.575 2.555 4.345 2.555 4.345 1.59 4.07 1.59  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.285 0.68 6.615 0.68 6.615 4.36 6.285 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 5.265 4.59 5.265 3.79 5.495 3.79 5.495 4.59 5.99 4.59 7.28 4.59 7.28 5.49 5.99 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 5.495 0.45 5.495 0.94 5.265 0.94 5.265 0.45 2.895 0.45 2.895 1.015 2.665 1.015 2.665 0.45 0.475 0.45 0.475 1.015 0.245 1.015 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.29 3.845 4.805 3.845 4.805 0.93 3.84 0.93 3.84 1.475 1.545 1.475 1.545 0.68 1.775 0.68 1.775 1.245 3.61 1.245 3.61 0.7 5.035 0.7 5.035 2.27 5.99 2.27 5.99 2.5 5.035 2.5 5.035 4.075 0.29 4.075  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.27 1.07 2.27 1.07 2.71 0.71 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 2.27 3.26 2.27 3.26 2.71 2.39 2.71  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 2.27 4.38 2.27 4.38 2.71 3.51 2.71  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 2.89 6.025 2.89 6.025 0.68 6.255 0.68 6.255 4.36 5.75 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 4.675 4.59 4.675 3.55 4.905 3.55 4.905 4.59 5.625 4.59 7.045 4.59 7.045 3.55 7.275 3.55 7.275 4.59 7.84 4.59 7.84 5.49 5.625 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 7.375 0.45 7.375 1.49 7.145 1.49 7.145 0.45 4.955 0.45 4.955 1.02 4.725 1.02 4.725 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 3.09 4.61 3.09 4.61 1.48 1.365 1.48 1.365 0.68 1.595 0.68 1.595 1.25 3.605 1.25 3.605 0.68 3.835 0.68 3.835 1.25 4.84 1.25 4.84 2.215 5.625 2.215 5.625 2.555 4.84 2.555 4.84 3.32 0.575 3.32 0.575 4.36 0.345 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.035 2.215 4.33 2.215 4.33 2.71 4.035 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.06 2.27 3.67 2.27 3.67 2.94 4.63 2.94 4.63 2.215 6.565 2.215 6.565 2.71 4.86 2.71 4.86 3.17 3.44 3.17 3.44 2.5 3.06 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.755 7.13 1.755 7.13 2.27 7.74 2.27 7.74 2.5 6.87 2.5 6.87 1.985 2.28 1.985 2.28 2.5 1.94 2.5  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.27 1.21 2.27 1.21 2.89 3.21 2.89 3.21 3.4 7.97 3.4 7.97 2.27 8.86 2.27 8.86 2.5 8.2 2.5 8.2 3.63 0.87 3.63  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5505 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.17 3.295 11.05 3.295 11.28 3.295 11.28 1.95 10.505 1.95 10.505 0.68 10.735 0.68 10.735 1.72 12.745 1.72 12.745 0.68 12.975 0.68 12.975 1.95 11.835 1.95 11.835 3.295 12.875 3.295 12.875 4.36 12.645 4.36 12.645 3.525 11.05 3.525 10.735 3.525 10.735 4.36 10.17 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.755 0.575 3.755 0.575 4.59 9.46 4.59 9.46 4.275 9.69 4.275 9.69 4.59 11.05 4.59 11.575 4.59 11.575 3.755 11.805 3.755 11.805 4.59 13.765 4.59 13.765 3.755 13.995 3.755 13.995 4.59 14.56 4.59 14.56 5.49 11.05 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 14.095 0.45 14.095 1.49 13.865 1.49 13.865 0.45 11.855 0.45 11.855 1.49 11.625 1.49 11.625 0.45 9.435 0.45 9.435 1.02 9.205 1.02 9.205 0.45 7.195 0.45 7.195 1.02 6.965 1.02 6.965 0.45 4.955 0.45 4.955 1.02 4.725 1.02 4.725 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.72 3.86 9.09 3.86 9.09 1.48 1.365 1.48 1.365 0.68 1.595 0.68 1.595 1.25 3.605 1.25 3.605 0.68 3.835 0.68 3.835 1.25 5.845 1.25 5.845 0.68 6.075 0.68 6.075 1.25 8.085 1.25 8.085 0.68 8.315 0.68 8.315 1.25 9.32 1.25 9.32 2.27 11.05 2.27 11.05 2.5 9.32 2.5 9.32 4.09 4.72 4.09  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.21 4.89 1.21 4.89 2.52 4.63 2.52  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.41 1.77 0.41 2.18 0.915 2.18 0.915 2.71 0.15 2.71  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.77 1.53 1.77 1.53 2.18 2.02 2.18 2.02 2.71 1.27 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 1.77 6.835 1.77 6.835 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.19 1.21 19.445 1.21 19.445 0.79 19.725 0.79 19.725 3.69 19.495 3.69 19.495 2.71 19.19 2.71  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.44 1.545 3.44 1.545 4.59 2.775 4.59 5.03 4.59 5.03 3.965 5.37 3.965 5.37 4.59 7.18 4.59 7.18 3.995 7.52 3.995 7.52 4.59 9.845 4.59 10.285 4.59 12.595 4.59 12.595 3.44 12.825 3.44 12.825 4.59 14.375 4.59 17.025 4.59 17.025 3.595 17.255 3.595 17.255 4.59 17.93 4.59 18.955 4.59 20.515 4.59 20.515 3.88 20.745 3.88 20.745 4.59 21.28 4.59 21.28 5.49 18.955 5.49 17.93 5.49 14.375 5.49 10.285 5.49 9.845 5.49 2.775 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.795 0.45 20.795 1.6 20.565 1.6 20.565 0.45 17.615 0.45 17.615 0.72 17.385 0.72 17.385 0.45 13.15 0.45 13.15 0.505 12.81 0.505 12.81 0.45 7.79 0.45 7.79 0.51 7.45 0.51 7.45 0.45 5.79 0.45 5.79 0.51 5.45 0.51 5.45 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 2.98 2.545 2.98 2.545 1.535 0.245 1.535 0.245 0.79 0.475 0.79 0.475 1.305 2.775 1.305 2.775 3.21 0.525 3.21 0.525 4.25 0.295 4.25  ;
        POLYGON 6.03 2.935 6.26 2.935 6.26 3.045 8.125 3.045 8.125 1.54 6.165 1.54 6.165 1.2 8.355 1.2 8.355 3.275 6.03 3.275  ;
        POLYGON 3.325 0.74 9.795 0.74 9.795 1.48 9.565 1.48 9.565 0.97 3.555 0.97 3.555 1.13 3.325 1.13  ;
        POLYGON 3.125 3.44 3.355 3.44 3.355 3.505 9.845 3.505 9.845 3.845 9.615 3.845 9.615 3.735 3.355 3.735 3.355 4.25 3.125 4.25  ;
        POLYGON 8.705 1.22 9.075 1.22 9.075 2.18 10.285 2.18 10.285 2.52 8.935 2.52 8.935 3.26 8.705 3.26  ;
        POLYGON 10.685 1.36 10.915 1.36 10.915 1.72 13.665 1.72 13.665 2.52 13.435 2.52 13.435 1.95 10.915 1.95 10.915 4.25 10.685 4.25  ;
        POLYGON 12.205 2.18 12.435 2.18 12.435 2.75 14.145 2.75 14.145 1.36 14.375 1.36 14.375 4.25 14.015 4.25 14.015 2.98 12.205 2.98  ;
        POLYGON 11.365 0.68 11.595 0.68 11.595 0.735 16.065 0.735 16.065 2.905 15.725 2.905 15.725 1.02 11.365 1.02  ;
        POLYGON 15.265 1.36 15.495 1.36 15.495 3.135 17.59 3.135 17.59 2.235 17.93 2.235 17.93 3.365 15.495 3.365 15.495 4.25 15.265 4.25  ;
        POLYGON 18.225 2.29 18.725 2.29 18.725 1.545 16.97 1.545 16.97 2.465 16.63 2.465 16.63 1.315 18.955 1.315 18.955 2.52 18.455 2.52 18.455 4.25 18.225 4.25  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 22.4 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.225 4.835 2.225 4.835 2.71 4.07 2.71  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.41 1.77 0.41 2.225 1.015 2.225 1.015 2.71 0.15 2.71  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.135 1.77 2.135 2.71 1.83 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 1.77 7.69 1.77 7.69 2.71 7.43 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.70205 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.79 0.845 21.13 0.845 21.13 4.25 20.79 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.44 1.595 3.44 1.595 4.59 2.895 4.59 5.235 4.59 5.235 3.905 5.465 3.905 5.465 4.59 7.83 4.59 7.83 3.905 8.17 3.905 8.17 4.59 10.685 4.59 11.125 4.59 13.235 4.59 13.235 3.44 13.465 3.44 13.465 4.59 14.485 4.59 17.645 4.59 17.645 3.6 17.875 3.6 17.875 4.59 18.37 4.59 19.41 4.59 19.735 4.59 19.735 3.88 19.965 3.88 19.965 4.59 21.81 4.59 21.81 3.88 22.04 3.88 22.04 4.59 22.4 4.59 22.4 5.49 19.41 5.49 18.37 5.49 14.485 5.49 11.125 5.49 10.685 5.49 2.895 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 22.4 -0.45 22.4 0.45 22.155 0.45 22.155 1.165 21.925 1.165 21.925 0.45 19.915 0.45 19.915 1.6 19.685 1.6 19.685 0.45 17.975 0.45 17.975 1.59 17.745 1.59 17.745 0.45 13.1 0.45 13.1 0.62 12.87 0.62 12.87 0.45 7.795 0.45 7.795 0.62 7.565 0.62 7.565 0.45 5.735 0.45 5.735 0.62 5.505 0.62 5.505 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.98 2.665 2.98 2.665 1.54 0.245 1.54 0.245 0.79 0.475 0.79 0.475 1.31 2.895 1.31 2.895 3.21 0.575 3.21 0.575 4.25 0.345 4.25  ;
        POLYGON 6.865 2.875 7.095 2.875 7.095 2.985 8.325 2.985 8.325 1.54 6.455 1.54 6.455 1.65 6.225 1.65 6.225 1.31 8.555 1.31 8.555 3.215 6.865 3.215  ;
        POLYGON 3.325 0.79 3.555 0.79 3.555 0.85 9.855 0.85 9.855 1.43 9.625 1.43 9.625 1.08 3.555 1.08 3.555 1.13 3.325 1.13  ;
        POLYGON 3.375 3.44 3.605 3.44 3.605 4.02 4.775 4.02 4.775 3.445 10.685 3.445 10.685 3.785 10.455 3.785 10.455 3.675 5.005 3.675 5.005 4.25 3.375 4.25  ;
        POLYGON 8.905 1.31 9.135 1.31 9.135 2.225 11.125 2.225 11.125 2.565 9.135 2.565 9.135 3.215 8.905 3.215  ;
        POLYGON 10.745 1.31 11.705 1.31 11.705 1.765 13.755 1.765 13.755 2.565 13.525 2.565 13.525 1.995 11.705 1.995 11.705 4.25 11.475 4.25 11.475 1.65 10.745 1.65  ;
        POLYGON 12.795 2.225 13.025 2.225 13.025 2.795 14.205 2.795 14.205 1.31 14.485 1.31 14.485 4.25 14.255 4.25 14.255 3.025 12.795 3.025  ;
        POLYGON 11.37 0.685 11.71 0.685 11.71 0.85 14.73 0.85 14.73 0.685 16.015 0.685 16.015 2.91 15.785 2.91 15.785 1.08 11.37 1.08  ;
        POLYGON 15.325 1.31 15.555 1.31 15.555 3.14 17.665 3.14 17.665 2.28 18.37 2.28 18.37 2.51 17.895 2.51 17.895 3.37 15.555 3.37 15.555 4.25 15.325 4.25  ;
        POLYGON 17.205 1.82 18.865 1.82 18.865 0.79 19.095 0.79 19.095 2.225 19.41 2.225 19.41 2.565 18.895 2.565 18.895 4.25 18.665 4.25 18.665 2.05 17.435 2.05 17.435 2.565 17.205 2.565  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.64 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.03 4.835 2.03 4.835 2.37 4.33 2.37 4.33 2.71 4.07 2.71  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.415 1.77 0.415 2.71 0.15 2.71  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.03 2.035 2.03 2.035 2.37 0.97 2.37 0.97 2.71 0.71 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 1.77 5.625 1.77 5.625 2.71 5.19 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.46815 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.705 0.845 20.935 0.845 20.935 1.92 22.55 1.92 22.55 1.21 22.945 1.21 22.945 0.845 23.175 0.845 23.175 1.655 22.81 1.655 22.81 2.15 20.935 2.15 20.935 3.415 23.035 3.415 23.035 4.25 22.805 4.25 22.805 3.645 20.985 3.645 20.985 4.25 20.705 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.465 4.59 10.52 4.59 11.095 4.59 13.085 4.59 13.085 3.44 13.315 3.44 13.315 4.59 14.435 4.59 17.645 4.59 17.645 3.55 17.875 3.55 17.875 4.59 18.44 4.59 19.735 4.59 19.735 3.875 19.965 3.875 19.965 4.59 20.255 4.59 21.775 4.59 21.775 3.875 22.005 3.875 22.005 4.59 23.93 4.59 23.93 3.875 24.16 3.875 24.16 4.59 24.64 4.59 24.64 5.49 20.255 5.49 18.44 5.49 14.435 5.49 11.095 5.49 10.52 5.49 3.055 5.49 0 5.49 0 4.59 1.645 4.59 1.645 3.44 1.875 3.44 1.875 4.59 3.055 4.59 5.235 4.59 5.235 3.905 8.17 3.905 8.17 4.135 5.465 4.135  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 24.64 -0.45 24.64 0.45 24.295 0.45 24.295 1.165 24.065 1.165 24.065 0.45 22.055 0.45 22.055 1.165 21.825 1.165 21.825 0.45 19.815 0.45 19.815 1.6 19.585 1.6 19.585 0.45 17.975 0.45 17.975 1.395 17.745 1.395 17.745 0.45 13.15 0.45 13.15 0.625 12.92 0.625 12.92 0.45 7.795 0.45 7.795 0.625 7.565 0.625 7.565 0.45 5.735 0.45 5.735 0.625 5.505 0.625 5.505 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.625 2.98 2.825 2.98 2.825 1.535 0.245 1.535 0.245 0.79 0.475 0.79 0.475 1.305 3.055 1.305 3.055 3.21 0.855 3.21 0.855 4.25 0.625 4.25  ;
        POLYGON 6.865 2.875 8.225 2.875 8.225 1.655 6.225 1.655 6.225 1.315 8.455 1.315 8.455 3.215 6.865 3.215  ;
        POLYGON 3.325 0.79 3.555 0.79 3.555 0.855 9.855 0.855 9.855 1.435 9.625 1.435 9.625 1.085 3.555 1.085 3.555 1.13 3.325 1.13  ;
        POLYGON 3.405 3.44 3.635 3.44 3.635 3.445 10.52 3.445 10.52 3.785 10.29 3.785 10.29 3.675 3.635 3.675 3.635 4.25 3.405 4.25  ;
        POLYGON 8.905 1.315 9.135 1.315 9.135 2.03 11.095 2.03 11.095 2.37 9.135 2.37 9.135 3.215 8.905 3.215  ;
        POLYGON 10.745 1.315 11.54 1.315 11.54 1.57 13.755 1.57 13.755 2.37 13.525 2.37 13.525 1.8 11.555 1.8 11.555 4.25 11.325 4.25 11.325 1.655 10.745 1.655  ;
        POLYGON 12.645 2.03 12.875 2.03 12.875 2.6 14.205 2.6 14.205 1.315 14.435 1.315 14.435 4.25 14.205 4.25 14.205 2.83 12.645 2.83  ;
        POLYGON 11.37 0.69 11.71 0.69 11.71 0.855 14.73 0.855 14.73 0.69 16.125 0.69 16.125 2.86 15.785 2.86 15.785 1.085 11.37 1.085  ;
        POLYGON 15.325 1.315 15.555 1.315 15.555 3.09 17.665 3.09 17.665 2.085 18.44 2.085 18.44 2.315 17.895 2.315 17.895 3.32 15.555 3.32 15.555 4.25 15.325 4.25  ;
        POLYGON 17.205 1.625 18.865 1.625 18.865 0.79 19.095 0.79 19.095 2.03 20.255 2.03 20.255 2.37 18.965 2.37 18.965 4.25 18.735 4.25 18.735 1.855 17.435 1.855 17.435 2.37 17.205 2.37  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 22.96 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 2.33 4.33 2.33 4.33 2.71 3.51 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.63 1.77 18.89 1.77 18.89 2.71 18.63 2.71  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.33 0.97 2.33 0.97 2.71 0.15 2.71  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.33 2.09 2.33 2.09 2.71 1.27 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.33 7.13 2.33 7.13 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.87 0.845 21.33 0.845 21.33 4.25 20.87 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.44 1.545 3.44 1.545 4.59 5.085 4.59 5.085 3.44 5.315 3.44 5.315 4.59 7.18 4.59 7.18 4.03 7.52 4.03 7.52 4.59 9.38 4.59 9.82 4.59 12.155 4.59 12.155 3.91 12.385 3.91 12.385 4.59 13.405 4.59 13.955 4.59 13.955 3.44 14.185 3.44 14.185 4.59 14.31 4.59 15.205 4.59 18.2 4.59 18.2 3.91 18.43 3.91 18.43 4.59 19.91 4.59 20.24 4.59 20.24 3.44 20.47 3.44 20.47 4.59 20.63 4.59 22.12 4.59 22.12 3.44 22.35 3.44 22.35 4.59 22.96 4.59 22.96 5.49 20.63 5.49 19.91 5.49 15.205 5.49 14.31 5.49 13.405 5.49 9.82 5.49 9.38 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 22.96 -0.45 22.96 0.45 22.4 0.45 22.4 1.655 22.17 1.655 22.17 0.45 18.43 0.45 18.43 1.275 18.2 1.275 18.2 0.45 13.495 0.45 13.495 1.44 13.265 1.44 13.265 0.45 7.515 0.45 7.515 1.18 7.285 1.18 7.285 0.45 5.68 0.45 5.68 0.53 5.45 0.53 5.45 0.45 1.595 0.45 1.595 1.285 1.365 1.285 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 2.98 2.545 2.98 2.545 2.1 0.245 2.1 0.245 0.945 0.475 0.945 0.475 1.87 4.835 1.87 4.835 2.635 4.605 2.635 4.605 2.1 2.775 2.1 2.775 3.21 0.525 3.21 0.525 4.25 0.295 4.25  ;
        POLYGON 6.16 3.01 7.725 3.01 7.725 2.1 6.165 2.1 6.165 1.21 6.395 1.21 6.395 1.87 7.955 1.87 7.955 3.24 6.16 3.24  ;
        POLYGON 3.325 0.76 6.025 0.76 6.025 0.75 6.855 0.75 6.855 1.41 7.945 1.41 7.945 0.68 9.355 0.68 9.355 1.275 9.125 1.275 9.125 0.91 8.175 0.91 8.175 1.64 6.625 1.64 6.625 0.98 6.095 0.98 6.095 0.99 3.555 0.99 3.555 1.285 3.325 1.285  ;
        POLYGON 3.325 2.98 5.775 2.98 5.775 3.525 9.38 3.525 9.38 3.755 5.545 3.755 5.545 3.21 3.555 3.21 3.555 4.25 3.325 4.25  ;
        POLYGON 8.305 2.39 8.405 2.39 8.405 1.14 8.635 1.14 8.635 2.35 9.82 2.35 9.82 2.58 8.535 2.58 8.535 3.295 8.305 3.295  ;
        POLYGON 11.135 3.44 13.405 3.44 13.405 4.25 13.175 4.25 13.175 3.67 11.365 3.67 11.365 4.25 11.135 4.25  ;
        POLYGON 10.115 0.945 10.475 0.945 10.475 2.865 13.97 2.865 13.97 2.59 14.31 2.59 14.31 3.095 10.345 3.095 10.345 4.25 10.115 4.25  ;
        POLYGON 11.765 2.13 14.605 2.13 14.605 1.155 14.835 1.155 14.835 2.205 15.205 2.205 15.205 4.25 14.975 4.25 14.975 2.435 14.665 2.435 14.665 2.36 11.995 2.36 11.995 2.635 11.765 2.635  ;
        POLYGON 10.825 1.67 14.145 1.67 14.145 0.695 16.83 0.695 16.83 3.15 16.6 3.15 16.6 0.925 15.295 0.925 15.295 1.955 15.065 1.955 15.065 0.925 14.375 0.925 14.375 1.9 11.055 1.9 11.055 2.635 10.825 2.635  ;
        POLYGON 17.08 1.155 17.41 1.155 17.41 3.78 17.08 3.78  ;
        POLYGON 15.67 1.21 16.225 1.21 16.225 4.02 17.74 4.02 17.74 3.45 18.89 3.45 18.89 4.01 19.68 4.01 19.68 2.295 19.91 2.295 19.91 4.24 18.66 4.24 18.66 3.68 17.97 3.68 17.97 4.25 15.995 4.25 15.995 1.44 15.67 1.44  ;
        POLYGON 17.76 2.295 17.99 2.295 17.99 2.94 19.22 2.94 19.22 1.835 20.24 1.835 20.24 0.945 20.63 0.945 20.63 2.635 20.4 2.635 20.4 2.065 19.45 2.065 19.45 3.78 19.22 3.78 19.22 3.17 17.76 3.17  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 2.33 3.995 2.33 3.995 3.27 3.51 3.27  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.144 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.07 2.89 18.61 2.89 18.61 1.77 18.89 1.77 18.89 3.27 18.07 3.27  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.33 1.53 2.33 1.53 2.735 0.71 2.735  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 1.83 2.15 1.83 2.15 2.75 1.77 2.75  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.33 7.13 2.33 7.13 2.735 6.31 2.735  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6746 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.895 0.84 22.25 0.84 22.25 4.25 21.895 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.44 1.595 3.44 1.595 4.59 5.085 4.59 5.085 3.44 5.315 3.44 5.315 4.59 7.175 4.59 7.175 3.94 7.515 3.94 7.515 4.59 9.2 4.59 9.695 4.59 12.03 4.59 12.03 3.44 12.26 3.44 12.26 4.59 13.28 4.59 13.77 4.59 13.77 3.44 13.955 3.44 14 3.44 14 4.59 15.02 4.59 18.07 4.59 18.07 4.48 18.3 4.48 18.3 4.59 20 4.59 20.33 4.59 20.33 3.44 20.56 3.44 20.56 4.59 20.585 4.59 22.915 4.59 22.915 3.44 23.145 3.44 23.145 4.59 23.52 4.59 23.52 5.49 20.585 5.49 20 5.49 15.02 5.49 13.955 5.49 13.28 5.49 9.695 5.49 9.2 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 23.275 0.45 23.275 1.16 23.045 1.16 23.045 0.45 21.035 0.45 21.035 1.16 20.805 1.16 20.805 0.45 18.08 0.45 18.08 1.325 17.85 1.325 17.85 0.45 13.36 0.45 13.36 1.325 13.13 1.325 13.13 0.45 7.56 0.45 7.56 1.18 7.33 1.18 7.33 0.45 5.735 0.45 5.735 0.605 5.505 0.605 5.505 0.45 1.595 0.45 1.595 1.14 1.365 1.14 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.98 2.545 2.98 2.545 1.6 0.245 1.6 0.245 0.8 0.475 0.8 0.475 1.37 4.99 1.37 4.99 2.735 4.65 2.735 4.65 1.6 2.775 1.6 2.775 3.21 0.575 3.21 0.575 4.25 0.345 4.25  ;
        POLYGON 6.155 2.965 7.36 2.965 7.36 2.1 6.21 2.1 6.21 1.27 6.44 1.27 6.44 1.87 7.59 1.87 7.59 2.505 7.955 2.505 7.955 2.735 7.59 2.735 7.59 3.195 6.155 3.195  ;
        POLYGON 3.125 3.44 3.355 3.44 3.355 4.02 4.625 4.02 4.625 2.98 5.775 2.98 5.775 3.48 8.97 3.48 8.97 3.44 9.2 3.44 9.2 4.25 8.97 4.25 8.97 3.71 5.545 3.71 5.545 3.21 4.855 3.21 4.855 4.25 3.125 4.25  ;
        POLYGON 3.27 0.835 6 0.835 6 0.81 6.9 0.81 6.9 1.41 7.99 1.41 7.99 0.755 9.42 0.755 9.42 1.325 9.19 1.325 9.19 0.985 8.22 0.985 8.22 1.64 6.67 1.64 6.67 1.04 6.105 1.04 6.105 1.065 3.61 1.065 3.61 1.085 3.27 1.085  ;
        POLYGON 8.25 2.52 8.45 2.52 8.45 1.215 8.68 1.215 8.68 2.505 9.695 2.505 9.695 2.735 8.535 2.735 8.535 3.25 8.25 3.25  ;
        POLYGON 11.01 2.98 13.28 2.98 13.28 4.25 13.05 4.25 13.05 3.21 11.24 3.21 11.24 4.25 11.01 4.25  ;
        POLYGON 9.99 2.685 10.31 2.685 10.31 0.985 10.54 0.985 10.54 2.505 13.955 2.505 13.955 2.735 10.535 2.735 10.535 2.915 10.22 2.915 10.22 4.25 9.99 4.25  ;
        POLYGON 11.535 2.045 14.25 2.045 14.25 1.215 14.48 1.215 14.48 3.02 15.02 3.02 15.02 4.25 14.79 4.25 14.79 3.25 14.25 3.25 14.25 2.275 11.535 2.275  ;
        POLYGON 10.835 1.585 13.79 1.585 13.79 0.755 16.5 0.755 16.5 2.79 16.27 2.79 16.27 0.985 15.02 0.985 15.02 2.79 14.79 2.79 14.79 0.985 14.02 0.985 14.02 1.815 11.175 1.815 11.175 1.96 10.835 1.96  ;
        POLYGON 16.73 1.215 17.06 1.215 17.06 3.78 16.73 3.78  ;
        POLYGON 15.39 1.215 16.04 1.215 16.04 4.02 19.77 4.02 19.77 2.525 20 2.525 20 4.25 15.81 4.25 15.81 1.555 15.39 1.555  ;
        POLYGON 17.41 2.45 17.64 2.45 17.64 3.55 19.31 3.55 19.31 1.985 19.99 1.985 19.99 0.8 20.22 0.8 20.22 1.985 20.585 1.985 20.585 2.215 19.54 2.215 19.54 3.78 17.41 3.78  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 26.32 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 2.33 4.49 2.33 4.49 2.735 3.51 2.735  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.144 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.63 1.77 18.89 1.77 18.89 2.79 18.63 2.79  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.175 1.77 1.175 2.735 0.71 2.735  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.53 1.77 2.53 2.735 1.83 2.735  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.87 1.77 7.4 1.77 7.4 2.735 6.87 2.735  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 22.425 0.84 22.655 0.84 22.655 1.39 24.23 1.39 24.23 1.21 24.665 1.21 24.665 0.84 24.895 0.84 24.895 4.25 24.23 4.25 24.23 1.62 22.655 1.62 22.655 4.25 22.425 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.51 4.59 1.51 3.44 1.74 3.44 1.74 4.59 5.525 4.59 5.525 3.44 5.755 3.44 5.755 4.59 7.64 4.59 7.64 3.94 7.98 3.94 7.98 4.59 9.995 4.59 10.49 4.59 12.825 4.59 12.825 3.45 13.055 3.45 13.055 4.59 14.075 4.59 14.585 4.59 14.585 3.44 14.77 3.44 14.815 3.44 14.815 4.59 15.835 4.59 18.885 4.59 18.885 4.35 19.115 4.35 19.115 4.59 20.595 4.59 20.925 4.59 20.925 3.44 21.085 3.44 21.155 3.44 21.155 4.59 23.495 4.59 23.495 3.44 23.725 3.44 23.725 4.59 25.645 4.59 25.645 3.44 25.875 3.44 25.875 4.59 26.32 4.59 26.32 5.49 21.085 5.49 20.595 5.49 15.835 5.49 14.77 5.49 14.075 5.49 10.49 5.49 9.995 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 26.32 -0.45 26.32 0.45 26.015 0.45 26.015 1.16 25.785 1.16 25.785 0.45 23.775 0.45 23.775 1.16 23.545 1.16 23.545 0.45 21.535 0.45 21.535 1.16 21.305 1.16 21.305 0.45 18.675 0.45 18.675 1.38 18.445 1.38 18.445 0.45 14.175 0.45 14.175 1.38 13.945 1.38 13.945 0.45 8.195 0.45 8.195 0.62 7.965 0.62 7.965 0.45 6.175 0.45 6.175 0.645 5.945 0.645 5.945 0.45 1.815 0.45 1.815 1.08 1.585 1.08 1.585 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.49 2.965 2.985 2.965 2.985 1.54 0.245 1.54 0.245 1.005 0.475 1.005 0.475 1.31 3.215 1.31 3.215 1.87 5.375 1.87 5.375 2.75 5.145 2.75 5.145 2.1 3.215 2.1 3.215 3.195 0.72 3.195 0.72 4.25 0.49 4.25  ;
        POLYGON 6.62 2.965 7.63 2.965 7.63 2.505 8.19 2.505 8.19 1.54 6.57 1.54 6.57 1.31 8.42 1.31 8.42 2.735 7.86 2.735 7.86 3.195 6.62 3.195  ;
        POLYGON 3.765 2.98 6.215 2.98 6.215 3.48 9.765 3.48 9.765 3.44 9.995 3.44 9.995 4.25 9.765 4.25 9.765 3.71 5.985 3.71 5.985 3.21 3.995 3.21 3.995 4.25 3.765 4.25  ;
        POLYGON 3.765 0.875 6.36 0.875 6.36 0.85 8.855 0.85 8.855 0.735 10.255 0.735 10.255 1.38 10.025 1.38 10.025 0.965 9.08 0.965 9.08 1.08 6.465 1.08 6.465 1.105 3.995 1.105 3.995 1.345 3.765 1.345  ;
        POLYGON 8.715 2.505 9.305 2.505 9.305 1.195 9.535 1.195 9.535 2.505 10.49 2.505 10.49 2.735 8.945 2.735 8.945 3.25 8.715 3.25  ;
        POLYGON 11.805 2.99 14.075 2.99 14.075 4.25 13.845 4.25 13.845 3.22 12.035 3.22 12.035 4.25 11.805 4.25  ;
        POLYGON 10.785 2.71 11.145 2.71 11.145 1.07 11.375 1.07 11.375 2.53 14.77 2.53 14.77 2.76 11.37 2.76 11.37 2.94 11.015 2.94 11.015 4.25 10.785 4.25  ;
        POLYGON 12.37 2.07 15.065 2.07 15.065 1.27 15.295 1.27 15.295 3.02 15.835 3.02 15.835 4.25 15.605 4.25 15.605 3.25 15.065 3.25 15.065 2.3 12.37 2.3  ;
        POLYGON 11.67 1.61 14.605 1.61 14.605 0.81 17.095 0.81 17.095 1.84 17.295 1.84 17.295 2.79 17.065 2.79 17.065 2.07 16.865 2.07 16.865 1.04 15.835 1.04 15.835 2.79 15.605 2.79 15.605 1.04 14.835 1.04 14.835 1.84 12.01 1.84 12.01 2.015 11.67 2.015  ;
        POLYGON 17.325 1.27 17.755 1.27 17.755 3.44 17.875 3.44 17.875 3.78 17.525 3.78 17.525 1.61 17.325 1.61  ;
        POLYGON 16.185 1.27 16.415 1.27 16.415 2.885 16.855 2.885 16.855 4.02 18.4 4.02 18.4 3.89 19.375 3.89 19.375 3.93 20.365 3.93 20.365 2.855 20.345 2.855 20.345 2.515 20.595 2.515 20.595 4.16 19.245 4.16 19.245 4.12 18.68 4.12 18.68 4.245 18.45 4.245 18.45 4.25 16.625 4.25 16.625 3.115 16.185 3.115  ;
        POLYGON 18.005 2.45 18.235 2.45 18.235 3.02 19.885 3.02 19.885 1.985 20.585 1.985 20.585 0.8 20.815 0.8 20.815 1.985 21.085 1.985 21.085 2.215 20.115 2.215 20.115 3.155 20.135 3.155 20.135 3.7 19.905 3.7 19.905 3.25 18.005 3.25  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 25.76 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.21 1.77 3.21 2.2 4.075 2.2 4.075 2.43 3.21 2.43 3.21 2.71 2.95 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.43 1.77 21.795 1.77 21.795 2.71 21.43 2.71  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.41 1.77 0.41 2.145 0.94 2.145 0.94 2.71 0.15 2.71  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.745 1.77 20.01 1.77 20.01 2.71 19.745 2.71  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.71 1.83 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.33 7.13 2.33 7.13 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 24.775 2.33 25.285 2.33 25.285 0.845 25.515 0.845 25.515 2.56 25.05 2.56 25.05 4.075 24.775 4.075  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.34 4.59 1.34 3.435 1.57 3.435 1.57 4.59 5.11 4.59 5.11 3.905 5.34 3.905 5.34 4.59 7.03 4.59 7.03 4.005 7.37 4.005 7.37 4.59 9.075 4.59 9.515 4.59 12.125 4.59 12.125 4.33 12.355 4.33 12.355 4.59 15.245 4.59 15.245 4.505 15.475 4.505 15.475 4.59 17.21 4.59 19.275 4.59 19.275 4.07 19.505 4.07 19.505 4.59 21.48 4.59 21.48 4.265 21.82 4.265 21.82 4.59 23.245 4.59 23.575 4.59 23.575 3.74 23.805 3.74 23.805 4.59 24.425 4.59 25.76 4.59 25.76 5.49 24.425 5.49 23.245 5.49 17.21 5.49 9.515 5.49 9.075 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 25.76 -0.45 25.76 0.45 24.395 0.45 24.395 1.6 24.165 1.6 24.165 0.45 21.31 0.45 21.31 1.08 20.97 1.08 20.97 0.45 13.655 0.45 13.655 1.425 13.425 1.425 13.425 0.45 7.615 0.45 7.615 1.135 7.385 1.135 7.385 0.45 5.76 0.45 5.76 0.535 5.53 0.535 5.53 0.45 1.675 0.45 1.675 1.08 1.335 1.08 1.335 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.32 2.94 2.49 2.94 2.49 1.54 0.27 1.54 0.27 0.795 0.5 0.795 0.5 1.31 2.72 1.31 2.72 2.94 4.73 2.94 4.73 2.145 4.96 2.145 4.96 3.17 0.55 3.17 0.55 4.075 0.32 4.075  ;
        POLYGON 6.065 2.94 7.525 2.94 7.525 2.055 6.265 2.055 6.265 1.225 6.495 1.225 6.495 1.825 7.755 1.825 7.755 3.28 6.065 3.28  ;
        POLYGON 3.35 3.435 5.73 3.435 5.73 3.545 8.845 3.545 8.845 2.965 9.075 2.965 9.075 3.775 5.53 3.775 5.53 3.665 3.58 3.665 3.58 4.245 3.35 4.245  ;
        POLYGON 3.35 0.765 6.955 0.765 6.955 1.365 8.045 1.365 8.045 0.765 9.455 0.765 9.455 1.425 9.225 1.425 9.225 0.995 8.275 0.995 8.275 1.595 6.725 1.595 6.725 0.995 3.58 0.995 3.58 1.135 3.35 1.135  ;
        POLYGON 8.105 2.255 8.505 2.255 8.505 1.225 8.735 1.225 8.735 2.145 9.515 2.145 9.515 2.485 8.335 2.485 8.335 3.27 8.105 3.27  ;
        POLYGON 10.885 3.265 13.555 3.265 13.555 3.605 10.885 3.605  ;
        POLYGON 9.865 2.895 10.345 2.895 10.345 1.085 10.575 1.085 10.575 2.715 14.485 2.715 14.485 2.605 14.715 2.605 14.715 2.945 10.57 2.945 10.57 3.125 10.095 3.125 10.095 3.945 9.865 3.945  ;
        POLYGON 14.045 3.265 14.945 3.265 14.945 2.375 12.095 2.375 12.095 2.485 11.865 2.485 11.865 2.145 15.905 2.145 15.905 1.315 16.715 1.315 16.715 3.895 16.485 3.895 16.485 1.545 16.135 1.545 16.135 2.375 15.175 2.375 15.175 3.605 14.045 3.605  ;
        POLYGON 10.39 3.87 15.825 3.87 15.825 4.125 17.21 4.125 17.21 4.355 15.65 4.355 15.65 4.275 15.42 4.275 15.42 4.1 10.73 4.1 10.73 4.35 10.39 4.35  ;
        POLYGON 10.925 1.655 15.445 1.655 15.445 0.68 18.835 0.68 18.835 2.485 18.605 2.485 18.605 0.91 15.675 0.91 15.675 1.885 11.155 1.885 11.155 2.485 10.925 2.485  ;
        POLYGON 18.145 1.315 18.375 1.315 18.375 2.715 19.065 2.715 19.065 0.795 19.295 0.795 19.295 1.31 20.525 1.31 20.525 3.77 20.295 3.77 20.295 1.54 19.295 1.54 19.295 2.945 18.755 2.945 18.755 3.31 18.525 3.31 18.525 2.945 18.145 2.945  ;
        POLYGON 17.025 1.315 17.735 1.315 17.735 3.61 19.965 3.61 19.965 4 20.61 4 20.61 3.985 21.025 3.985 21.025 3.76 23.015 3.76 23.015 2.145 23.245 2.145 23.245 3.99 21.255 3.99 21.255 4.215 20.695 4.215 20.695 4.23 19.735 4.23 19.735 3.84 17.735 3.84 17.735 3.95 17.505 3.95 17.505 1.655 17.025 1.655  ;
        POLYGON 20.82 1.31 23.445 1.31 23.445 0.795 23.69 0.795 23.69 1.83 24.425 1.83 24.425 2.485 24.195 2.485 24.195 2.06 23.46 2.06 23.46 1.54 22.785 1.54 22.785 3.53 22.555 3.53 22.555 1.54 21.16 1.54 21.16 2.43 20.82 2.43  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 26.88 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 4.33 1.77 4.33 2.29 3.51 2.29  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.43 1.77 21.69 1.77 21.69 2.015 21.935 2.015 21.935 2.355 21.69 2.355 21.69 2.71 21.43 2.71  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.97 1.77 0.97 2.3 0.15 2.3  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.75 1.77 20.04 1.77 20.04 2.71 19.75 2.71  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.77 2.09 1.77 2.09 2.345 1.27 2.345  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.33 7.13 2.33 7.13 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 25.145 0.79 25.61 0.79 25.61 2.71 25.375 2.71 25.375 4.08 25.145 4.08  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.415 4.59 1.415 3.27 1.645 3.27 1.645 4.59 5.085 4.59 5.085 3.44 5.315 3.44 5.315 4.59 7.19 4.59 7.19 4.125 7.53 4.125 7.53 4.59 9.215 4.59 9.655 4.59 9.695 4.59 12.21 4.59 12.21 4.565 12.55 4.565 12.55 4.59 15.35 4.59 15.35 4.565 15.69 4.565 15.69 4.59 17.31 4.59 19.395 4.59 19.395 3.91 19.625 3.91 19.625 4.59 21.665 4.59 21.665 4.3 21.895 4.3 21.895 4.59 23.375 4.59 23.725 4.59 23.725 3.27 23.955 3.27 23.955 4.59 24.835 4.59 26.165 4.59 26.165 3.27 26.395 3.27 26.395 4.59 26.88 4.59 26.88 5.49 24.835 5.49 23.375 5.49 17.31 5.49 9.695 5.49 9.655 5.49 9.215 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 26.88 -0.45 26.88 0.45 26.635 0.45 26.635 1.6 26.405 1.6 26.405 0.45 24.395 0.45 24.395 1.6 24.165 1.6 24.165 0.45 21.31 0.45 21.31 1.08 20.97 1.08 20.97 0.45 13.775 0.45 13.775 1.48 13.545 1.48 13.545 0.45 7.775 0.45 7.775 1.08 7.545 1.08 7.545 0.45 5.735 0.45 5.735 1.08 5.505 1.08 5.505 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.395 2.575 2.595 2.575 2.595 1.54 0.245 1.54 0.245 0.79 0.475 0.79 0.475 1.31 2.825 1.31 2.825 2.52 4.605 2.52 4.605 2.015 4.835 2.015 4.835 2.75 2.745 2.75 2.745 2.805 0.625 2.805 0.625 4.08 0.395 4.08  ;
        POLYGON 6.225 3.095 7.36 3.095 7.36 2 6.425 2 6.425 1.17 6.655 1.17 6.655 1.77 8.215 1.77 8.215 2.11 7.59 2.11 7.59 3.435 6.225 3.435  ;
        POLYGON 3.325 2.98 5.775 2.98 5.775 3.665 8.985 3.665 8.985 3.085 9.215 3.085 9.215 3.895 5.545 3.895 5.545 3.21 3.555 3.21 3.555 4.08 3.325 4.08  ;
        POLYGON 8.265 2.335 8.665 2.335 8.665 1.17 8.895 1.17 8.895 2.225 9.655 2.225 9.655 2.565 8.495 2.565 8.495 3.435 8.265 3.435  ;
        POLYGON 3.325 0.79 3.555 0.79 3.555 1.31 5.965 1.31 5.965 0.71 7.115 0.71 7.115 1.31 8.205 1.31 8.205 0.71 9.695 0.71 9.695 1.48 9.465 1.48 9.465 0.94 8.435 0.94 8.435 1.54 6.885 1.54 6.885 0.94 6.195 0.94 6.195 1.54 3.325 1.54  ;
        POLYGON 11.025 3.27 13.675 3.27 13.675 3.61 11.025 3.61  ;
        POLYGON 10.005 2.74 10.585 2.74 10.585 1.37 10.815 1.37 10.815 2.74 14.535 2.74 14.535 3.08 14.305 3.08 14.305 2.97 10.235 2.97 10.235 3.93 10.005 3.93  ;
        POLYGON 14.165 3.535 15.905 3.535 15.905 2.51 12.005 2.51 12.005 2.17 15.905 2.17 15.905 1.37 16.135 1.37 16.135 3.645 16.585 3.645 16.585 3.065 16.815 3.065 16.815 3.875 14.165 3.875  ;
        POLYGON 10.53 4.105 17.31 4.105 17.31 4.335 10.53 4.335  ;
        POLYGON 11.165 1.71 15.445 1.71 15.445 0.68 18.835 0.68 18.835 2.355 18.605 2.355 18.605 1.02 15.675 1.02 15.675 1.94 11.395 1.94 11.395 2.355 11.165 2.355  ;
        POLYGON 18.145 1.37 18.375 1.37 18.375 2.585 19.065 2.585 19.065 1.025 19.295 1.025 19.295 1.31 20.63 1.31 20.63 3.27 20.645 3.27 20.645 3.61 20.4 3.61 20.4 1.54 19.295 1.54 19.295 2.815 18.855 2.815 18.855 3.305 18.625 3.305 18.625 2.815 18.145 2.815  ;
        POLYGON 17.025 1.37 17.255 1.37 17.255 2.74 17.835 2.74 17.835 3.535 19.035 3.535 19.035 3.45 20.085 3.45 20.085 3.84 23.145 3.84 23.145 2.415 23.375 2.415 23.375 4.07 19.855 4.07 19.855 3.68 19.215 3.68 19.215 3.765 17.605 3.765 17.605 2.97 17.025 2.97  ;
        POLYGON 20.86 1.31 23.445 1.31 23.445 0.845 23.675 0.845 23.675 1.965 24.835 1.965 24.835 2.355 24.605 2.355 24.605 2.195 23.445 2.195 23.445 1.54 22.915 1.54 22.915 3.61 22.685 3.61 22.685 1.54 21.2 1.54 21.2 2.3 20.86 2.3  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 29.12 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 3.77 1.77 3.77 2.71 3.51 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.43 2.215 21.69 2.215 21.69 3.27 21.43 3.27  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.27 0.97 2.27 0.97 2.71 0.15 2.71  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.13 2.95 19.655 2.95 19.655 2.74 20.01 2.74 20.01 3.27 19.13 3.27  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.27 2.09 2.27 2.09 2.71 1.27 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 2.89 6.28 2.89 6.28 2.53 6.57 2.53 6.57 3.27 5.75 3.27  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 24.85 2.89 25.25 2.89 25.25 0.845 25.48 0.845 25.48 2.89 27.49 2.89 27.49 0.845 27.72 0.845 27.72 3.12 26.73 3.12 26.73 3.44 27.12 3.44 27.12 4.25 26.47 4.25 26.47 3.12 25.08 3.12 25.08 4.25 24.85 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.44 1.495 3.44 1.495 4.59 4.95 4.59 4.95 4.56 5.29 4.56 5.29 4.59 6.885 4.59 6.885 4.56 7.225 4.56 7.225 4.59 9.13 4.59 9.57 4.59 9.61 4.59 12.12 4.59 12.12 4.51 12.35 4.51 12.35 4.59 15.32 4.59 15.32 4.51 15.55 4.51 15.55 4.59 17.355 4.59 19.39 4.59 19.39 3.985 19.62 3.985 19.62 4.59 21.595 4.59 21.595 4.375 21.935 4.375 21.935 4.59 23.36 4.59 23.71 4.59 23.71 3.44 23.94 3.44 23.94 4.59 24.8 4.59 25.87 4.59 25.87 3.44 26.1 3.44 26.1 4.59 27.91 4.59 27.91 3.44 28.14 3.44 28.14 4.59 29.12 4.59 29.12 5.49 24.8 5.49 23.36 5.49 17.355 5.49 9.61 5.49 9.57 5.49 9.13 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 29.12 -0.45 29.12 0.45 28.84 0.45 28.84 1.65 28.61 1.65 28.61 0.45 26.6 0.45 26.6 1.65 26.37 1.65 26.37 0.45 24.36 0.45 24.36 1.525 24.13 1.525 24.13 0.45 21.22 0.45 21.22 1.255 20.99 1.255 20.99 0.45 13.69 0.45 13.69 1.535 13.46 1.535 13.46 0.45 7.69 0.45 7.69 1.38 7.46 1.38 7.46 0.45 5.675 0.45 5.675 0.53 5.445 0.53 5.445 0.45 1.595 0.45 1.595 1.535 1.365 1.535 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.94 2.445 2.94 2.445 2.04 0.245 2.04 0.245 1.195 0.475 1.195 0.475 1.81 2.675 1.81 2.675 2.94 4.605 2.94 4.605 2.215 4.835 2.215 4.835 3.17 0.475 3.17 0.475 4.25 0.245 4.25  ;
        POLYGON 5.7 3.5 7.6 3.5 7.6 2.3 6.34 2.3 6.34 1.22 6.57 1.22 6.57 2.07 7.83 2.07 7.83 3.84 5.7 3.84  ;
        POLYGON 3.025 3.44 3.255 3.44 3.255 4.1 8.9 4.1 8.9 3.065 9.13 3.065 9.13 4.33 3.025 4.33  ;
        POLYGON 8.18 2.325 8.58 2.325 8.58 1.22 8.81 1.22 8.81 2.215 9.57 2.215 9.57 2.555 8.41 2.555 8.41 3.87 8.18 3.87  ;
        POLYGON 3.325 0.76 7.03 0.76 7.03 1.61 8.12 1.61 8.12 0.76 9.61 0.76 9.61 1.535 9.38 1.535 9.38 0.99 8.35 0.99 8.35 1.84 6.8 1.84 6.8 0.99 3.555 0.99 3.555 1.535 3.325 1.535  ;
        POLYGON 10.94 3.44 13.59 3.44 13.59 3.78 10.94 3.78  ;
        POLYGON 9.92 2.985 10.5 2.985 10.5 1.195 10.73 1.195 10.73 2.98 14.75 2.98 14.75 3.32 14.52 3.32 14.52 3.21 10.55 3.21 10.55 3.215 10.15 3.215 10.15 3.875 9.92 3.875  ;
        POLYGON 14.08 3.44 14.31 3.44 14.31 3.55 15.64 3.55 15.64 2.565 11.92 2.565 11.92 2.225 15.64 2.225 15.64 1.195 15.87 1.195 15.87 3.44 16.86 3.44 16.86 3.78 14.08 3.78  ;
        POLYGON 10.445 4.05 17.355 4.05 17.355 4.28 10.445 4.28  ;
        POLYGON 11.08 1.765 15.18 1.765 15.18 0.68 18.68 0.68 18.68 2.22 18.34 2.22 18.34 0.91 15.41 0.91 15.41 1.995 11.31 1.995 11.31 2.115 11.08 2.115  ;
        POLYGON 17.88 1.195 18.11 1.195 18.11 2.45 19.03 2.45 19.03 1.145 19.26 1.145 19.26 2.28 20.64 2.28 20.64 3.685 20.41 3.685 20.41 2.51 19.255 2.51 19.255 2.68 18.9 2.68 18.9 3.295 18.67 3.295 18.67 2.68 17.88 2.68  ;
        POLYGON 16.76 1.195 16.99 1.195 16.99 2.945 17.88 2.945 17.88 3.525 20.08 3.525 20.08 3.915 23.13 3.915 23.13 2.215 23.36 2.215 23.36 4.145 19.85 4.145 19.85 3.755 17.65 3.755 17.65 3.175 16.76 3.175  ;
        POLYGON 20.795 1.755 23.41 1.755 23.41 0.845 23.64 0.845 23.64 1.755 24.8 1.755 24.8 2.555 24.57 2.555 24.57 1.985 22.9 1.985 22.9 3.685 22.67 3.685 22.67 1.985 21.135 1.985 21.135 2.11 20.795 2.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.64 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 3.995 1.77 3.995 2.71 3.51 2.71  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.275 0.97 2.275 0.97 2.71 0.15 2.71  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.63 1.77 19.425 1.77 19.425 2.71 18.63 2.71  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.275 2.09 2.275 2.09 2.71 1.27 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.275 7.13 2.275 7.13 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.67 0.845 24.285 0.845 24.285 4.06 23.67 4.06  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.4 1.545 3.4 1.545 4.59 5.145 4.59 5.145 3.25 5.375 3.25 5.375 4.59 7.45 4.59 7.45 3.97 7.79 3.97 7.79 4.59 9.675 4.59 10.17 4.59 12.595 4.59 12.595 3.835 12.825 3.835 12.825 4.59 14.955 4.59 14.955 3.09 15.185 3.09 15.185 4.59 16.865 4.59 18.955 4.59 18.955 3.4 19.185 3.4 19.185 4.59 20.205 4.59 21.195 4.59 21.195 4.31 21.425 4.31 21.425 4.59 22.985 4.59 22.985 3.25 23.215 3.25 23.215 4.59 23.44 4.59 24.64 4.59 24.64 5.49 23.44 5.49 20.205 5.49 16.865 5.49 10.17 5.49 9.675 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 24.64 -0.45 24.64 0.45 23.165 0.45 23.165 1.165 22.935 1.165 22.935 0.45 21.105 0.45 21.105 0.61 20.875 0.61 20.875 0.45 12.98 0.45 12.98 0.625 12.64 0.625 12.64 0.45 7.785 0.45 7.785 1.14 7.555 1.14 7.555 0.45 5.685 0.45 5.685 0.63 5.455 0.63 5.455 0.45 1.595 0.45 1.595 1.45 1.365 1.45 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 2.94 2.545 2.94 2.545 2.045 0.245 2.045 0.245 1.11 0.475 1.11 0.475 1.815 2.775 1.815 2.775 2.94 4.225 2.94 4.225 1.73 4.835 1.73 4.835 2.07 4.455 2.07 4.455 3.17 0.525 3.17 0.525 4.06 0.295 4.06  ;
        POLYGON 6.485 2.94 7.445 2.94 7.445 2.06 7.215 2.06 7.215 2.045 6.435 2.045 6.435 1.14 6.665 1.14 6.665 1.815 7.3 1.815 7.3 1.83 7.675 1.83 7.675 2.275 8.28 2.275 8.28 2.505 7.675 2.505 7.675 3.28 6.485 3.28  ;
        POLYGON 3.325 0.86 5.985 0.86 5.985 0.68 7.125 0.68 7.125 1.355 7.47 1.355 7.47 1.37 8.015 1.37 8.015 0.68 9.625 0.68 9.625 1.135 9.395 1.135 9.395 0.91 8.245 0.91 8.245 1.6 7.385 1.6 7.385 1.585 6.895 1.585 6.895 0.91 6.21 0.91 6.21 1.09 3.555 1.09 3.555 1.45 3.325 1.45  ;
        POLYGON 3.325 3.4 4.685 3.4 4.685 2.79 5.835 2.79 5.835 3.51 9.445 3.51 9.445 2.93 9.675 2.93 9.675 3.74 5.605 3.74 5.605 3.02 4.915 3.02 4.915 3.63 3.555 3.63 3.555 4.21 3.325 4.21  ;
        POLYGON 8.575 1.14 8.905 1.14 8.905 2.275 10.17 2.275 10.17 2.505 8.805 2.505 8.805 3.235 8.575 3.235  ;
        POLYGON 10.515 1.025 10.745 1.025 10.745 2.055 13.64 2.055 13.64 2.285 10.745 2.285 10.745 3.73 10.515 3.73  ;
        POLYGON 11.195 0.855 15.44 0.855 15.44 0.68 15.78 0.68 15.78 1.085 11.425 1.085 11.425 1.825 11.195 1.825  ;
        POLYGON 11.88 2.515 13.935 2.515 13.935 1.315 15.285 1.315 15.285 1.68 16.425 1.68 16.425 3.73 16.195 3.73 16.195 1.91 15.055 1.91 15.055 1.545 14.165 1.545 14.165 3.26 13.935 3.26 13.935 2.745 11.88 2.745  ;
        POLYGON 11.095 3.375 13.225 3.375 13.225 3.49 14.495 3.49 14.495 2.63 15.965 2.63 15.965 4.02 16.865 4.02 16.865 4.36 15.735 4.36 15.735 2.86 14.725 2.86 14.725 3.72 13.025 3.72 13.025 3.605 11.325 3.605 11.325 4.36 11.095 4.36  ;
        POLYGON 18.4 2.94 20.205 2.94 20.205 3.95 19.975 3.95 19.975 3.17 18.465 3.17 18.465 3.9 18.17 3.9 18.17 1.48 17.295 1.48 17.295 1.14 18.985 1.14 18.985 1.48 18.4 1.48  ;
        POLYGON 16.175 0.68 19.425 0.68 19.425 0.84 21.865 0.84 21.865 2.56 21.635 2.56 21.635 1.07 19.205 1.07 19.205 0.91 17.065 0.91 17.065 1.71 17.445 1.71 17.445 3.9 17.215 3.9 17.215 1.94 16.835 1.94 16.835 0.91 16.405 0.91 16.405 1.45 16.175 1.45  ;
        POLYGON 20.555 2.22 20.785 2.22 20.785 2.79 22.215 2.79 22.215 1.11 22.445 1.11 22.445 2.22 23.44 2.22 23.44 2.56 22.445 2.56 22.445 4.1 22.215 4.1 22.215 3.02 20.555 3.02  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 25.2 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 4.07 1.77 4.07 2.71 3.51 2.71  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.32 1.53 2.32 1.53 2.71 0.71 2.71  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.63 1.21 18.89 1.21 18.89 2.265 19.11 2.265 19.11 2.605 18.63 2.605  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.32 2.65 2.32 2.65 2.71 1.83 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.865 2.32 7.69 2.32 7.69 2.71 6.865 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.605 0.845 23.93 0.845 23.93 4.05 23.605 4.05  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.44 4.59 1.44 3.4 1.67 3.4 1.67 4.59 5.16 4.59 5.16 3.76 5.39 3.76 5.39 4.59 7.36 4.59 7.36 3.86 7.59 3.86 7.59 4.59 9.48 4.59 9.975 4.59 12.28 4.59 12.28 3.56 12.51 3.56 12.51 4.59 14.54 4.59 14.54 3.56 14.77 3.56 14.77 4.59 16.33 4.59 18.44 4.59 18.44 3.295 18.67 3.295 18.67 4.59 19.69 4.59 20.48 4.59 20.48 3.24 20.71 3.24 20.71 4.59 22.585 4.59 22.585 3.24 22.815 3.24 22.815 4.59 23.255 4.59 24.625 4.59 24.625 3.24 24.855 3.24 24.855 4.59 25.2 4.59 25.2 5.49 23.255 5.49 19.69 5.49 16.33 5.49 9.975 5.49 9.48 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 25.2 -0.45 25.2 0.45 24.955 0.45 24.955 1.165 24.725 1.165 24.725 0.45 22.715 0.45 22.715 1.165 22.485 1.165 22.485 0.45 20.61 0.45 20.61 1.48 20.38 1.48 20.38 0.45 12.51 0.45 12.51 1.22 12.28 1.22 12.28 0.45 7.59 0.45 7.59 1.17 7.36 1.17 7.36 0.45 5.775 0.45 5.775 0.575 5.545 0.575 5.545 0.45 1.67 0.45 1.67 1.48 1.44 1.48 1.44 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.94 2.88 2.94 2.88 2.09 0.32 2.09 0.32 1.14 0.55 1.14 0.55 1.86 3.11 1.86 3.11 2.94 4.4 2.94 4.4 2.84 4.68 2.84 4.68 2.265 4.91 2.265 4.91 3.07 4.59 3.07 4.59 3.17 0.65 3.17 0.65 4.05 0.42 4.05  ;
        POLYGON 6.34 2.875 6.57 2.875 6.57 2.94 7.92 2.94 7.92 2.09 6.24 2.09 6.24 1.26 6.47 1.26 6.47 1.86 8.15 1.86 8.15 3.17 6.57 3.17 6.57 3.215 6.34 3.215  ;
        POLYGON 3.4 0.805 6.14 0.805 6.14 0.8 6.93 0.8 6.93 1.4 7.82 1.4 7.82 0.68 9.43 0.68 9.43 1.22 9.2 1.22 9.2 0.91 8.05 0.91 8.05 1.63 6.7 1.63 6.7 1.03 6.19 1.03 6.19 1.035 3.63 1.035 3.63 1.48 3.4 1.48  ;
        POLYGON 3.4 3.4 4.78 3.4 4.78 3.3 5.82 3.3 5.82 3.445 7.08 3.445 7.08 3.4 8.05 3.4 8.05 3.915 9.25 3.915 9.25 3.09 9.48 3.09 9.48 4.145 7.82 4.145 7.82 3.63 7.22 3.63 7.22 3.675 5.605 3.675 5.605 3.53 4.97 3.53 4.97 3.63 3.63 3.63 3.63 4.21 3.4 4.21  ;
        POLYGON 8.38 1.14 8.71 1.14 8.71 2.32 9.975 2.32 9.975 2.55 8.61 2.55 8.61 3.685 8.38 3.685  ;
        POLYGON 10.32 1.11 10.55 1.11 10.55 2.085 11.555 2.085 11.555 2.055 13.225 2.055 13.225 2.285 11.67 2.285 11.67 2.315 10.55 2.315 10.55 3.73 10.32 3.73  ;
        POLYGON 10.845 1.595 12.74 1.595 12.74 0.68 15.265 0.68 15.265 0.91 12.97 0.91 12.97 1.825 11.185 1.825 11.185 1.855 10.845 1.855  ;
        POLYGON 11.785 2.515 14.54 2.515 14.54 1.14 14.77 1.14 14.77 2.515 15.89 2.515 15.89 3.685 15.66 3.685 15.66 2.745 13.75 2.745 13.75 3.73 13.52 3.73 13.52 2.745 11.785 2.745  ;
        POLYGON 10.9 3.1 12.97 3.1 12.97 3.96 14.08 3.96 14.08 3.1 15.43 3.1 15.43 3.975 16.33 3.975 16.33 4.315 15.2 4.315 15.2 3.33 14.31 3.33 14.31 4.19 12.74 4.19 12.74 3.33 11.13 3.33 11.13 4.36 10.9 4.36  ;
        POLYGON 17.72 2.835 18.17 2.835 18.17 1.655 16.78 1.655 16.78 1.315 18.4 1.315 18.4 2.835 19.69 2.835 19.69 4.05 19.46 4.05 19.46 3.065 17.95 3.065 17.95 3.845 17.72 3.845  ;
        POLYGON 15.66 1.14 16.32 1.14 16.32 0.75 19.35 0.75 19.35 1.71 20.73 1.71 20.73 2.32 21.385 2.32 21.385 2.55 20.5 2.55 20.5 1.94 19.12 1.94 19.12 0.98 16.55 0.98 16.55 1.885 16.91 1.885 16.91 3.845 16.68 3.845 16.68 2.115 16.32 2.115 16.32 1.48 15.66 1.48  ;
        POLYGON 20.04 2.265 20.27 2.265 20.27 2.78 21.68 2.78 21.68 0.845 21.91 0.845 21.91 2.78 23.025 2.78 23.025 2.265 23.255 2.265 23.255 3.01 21.91 3.01 21.91 4.05 21.68 4.05 21.68 3.01 20.04 3.01  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 27.44 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 4.33 1.77 4.33 2.215 3.51 2.215  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.97 1.77 0.97 2.215 0.15 2.215  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.07 1.77 18.89 1.77 18.89 2.215 18.07 2.215  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.77 2.09 1.77 2.09 2.215 1.27 2.215  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 2.33 6.91 2.33 6.91 2.71 5.75 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.55965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.59 0.845 23.82 0.845 23.82 1.21 25.83 1.21 25.83 0.845 26.06 0.845 26.06 1.655 23.93 1.655 23.93 2.88 25.92 2.88 25.92 3.69 25.69 3.69 25.69 3.11 23.87 3.11 23.87 3.69 23.59 3.69  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.23 1.545 3.23 1.545 4.59 5.085 4.59 5.085 3.4 5.315 3.4 5.315 4.59 7.2 4.59 7.2 4.125 7.54 4.125 7.54 4.59 9.275 4.59 9.72 4.59 12.045 4.59 12.045 4.51 12.275 4.51 12.275 4.59 14.305 4.59 14.305 4.07 14.535 4.07 14.535 4.59 16.235 4.59 18.305 4.59 18.305 3.075 18.535 3.075 18.535 4.59 19.555 4.59 20.565 4.59 20.565 3.88 20.795 3.88 20.795 4.59 22.605 4.59 22.605 3.88 22.835 3.88 22.835 4.59 23.275 4.59 24.66 4.59 24.66 3.88 24.89 3.88 24.89 4.59 26.85 4.59 26.85 3.88 27.08 3.88 27.08 4.59 27.44 4.59 27.44 5.49 23.275 5.49 19.555 5.49 16.235 5.49 9.72 5.49 9.275 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 27.44 -0.45 27.44 0.45 27.18 0.45 27.18 1.655 26.95 1.655 26.95 0.45 24.94 0.45 24.94 0.98 24.71 0.98 24.71 0.45 22.7 0.45 22.7 1.655 22.47 1.655 22.47 0.45 20.46 0.45 20.46 1.265 20.23 1.265 20.23 0.45 12.455 0.45 12.455 1.12 12.225 1.12 12.225 0.45 7.535 0.45 7.535 1.18 7.305 1.18 7.305 0.45 5.735 0.45 5.735 0.53 5.505 0.53 5.505 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 2.455 2.545 2.455 2.545 1.54 0.245 1.54 0.245 0.925 0.475 0.925 0.475 1.31 2.775 1.31 2.775 2.455 4.605 2.455 4.605 1.93 4.835 1.93 4.835 2.685 0.525 2.685 0.525 4.04 0.295 4.04  ;
        POLYGON 6.235 3.095 7.14 3.095 7.14 2.1 6.185 2.1 6.185 1.27 6.415 1.27 6.415 1.87 7.98 1.87 7.98 2.215 7.37 2.215 7.37 3.435 6.235 3.435  ;
        POLYGON 3.325 2.94 5.775 2.94 5.775 3.665 9.045 3.665 9.045 3.065 9.275 3.065 9.275 3.895 5.545 3.895 5.545 3.17 3.555 3.17 3.555 4.04 3.325 4.04  ;
        POLYGON 3.325 0.76 6.875 0.76 6.875 1.41 7.965 1.41 7.965 0.76 9.375 0.76 9.375 1.12 9.145 1.12 9.145 0.99 8.195 0.99 8.195 1.64 6.645 1.64 6.645 0.99 3.555 0.99 3.555 1.13 3.325 1.13  ;
        POLYGON 8.275 3.095 8.425 3.095 8.425 1.22 8.655 1.22 8.655 1.985 9.72 1.985 9.72 2.215 8.655 2.215 8.655 3.435 8.275 3.435  ;
        POLYGON 10.065 0.925 10.495 0.925 10.495 1.985 13.17 1.985 13.17 2.215 10.295 2.215 10.295 3.875 10.065 3.875  ;
        POLYGON 10.79 1.525 12.685 1.525 12.685 0.68 15.13 0.68 15.13 0.91 12.915 0.91 12.915 1.755 10.79 1.755  ;
        POLYGON 11.33 2.445 14.405 2.445 14.405 1.315 14.635 1.315 14.635 2.445 15.775 2.445 15.775 3.38 15.545 3.38 15.545 2.675 13.515 2.675 13.515 3.77 13.285 3.77 13.285 2.675 11.33 2.675  ;
        POLYGON 10.59 4.05 13.745 4.05 13.745 3.095 13.975 3.095 13.975 3.61 16.005 3.61 16.005 3.095 16.235 3.095 16.235 4.36 16.005 4.36 16.005 3.84 13.975 3.84 13.975 4.28 10.59 4.28  ;
        POLYGON 17.815 2.615 19.555 2.615 19.555 3.715 19.325 3.715 19.325 2.845 17.815 2.845 17.815 3.9 17.585 3.9 17.585 1.5 16.645 1.5 16.645 1.16 18.32 1.16 18.32 1.5 17.815 1.5  ;
        POLYGON 15.525 1.085 16.185 1.085 16.185 0.7 19.35 0.7 19.35 1.985 21.055 1.985 21.055 2.215 19.12 2.215 19.12 0.93 16.415 0.93 16.415 1.73 16.795 1.73 16.795 3.9 16.565 3.9 16.565 1.96 16.185 1.96 16.185 1.425 15.525 1.425  ;
        POLYGON 19.905 2.445 21.35 2.445 21.35 0.845 21.58 0.845 21.58 2.42 23.275 2.42 23.275 2.76 21.815 2.76 21.815 3.69 21.585 3.69 21.585 2.785 19.905 2.785  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__tieh
  CLASS core gf180mcu_fd_sc_mcu9t5v0__tiehIGH ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__tieh 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.24 BY 5.04 ;
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.89 1.53 2.89 1.53 3.7 1.27 3.7  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.25 4.59 0.25 2.945 0.48 2.945 0.48 4.59 1.6 4.59 2.24 4.59 2.24 5.49 1.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.24 -0.45 2.24 0.45 0.48 0.45 0.48 1.355 0.25 1.355 0.25 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.875 1.83 1.37 1.83 1.37 1.315 1.6 1.315 1.6 2.06 0.875 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__tieh
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__tiel
  CLASS core gf180mcu_fd_sc_mcu9t5v0__tielOW ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__tiel 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.24 BY 5.04 ;
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.2904 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.215 1.21 1.595 1.21 1.595 1.59 1.215 1.59  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 2.945 0.575 2.945 0.575 4.59 1.595 4.59 2.24 4.59 2.24 5.49 1.595 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.24 -0.45 2.24 0.45 0.475 0.45 0.475 1.355 0.245 1.355 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.87 2.47 1.595 2.47 1.595 3.685 1.365 3.685 1.365 2.7 0.87 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__tiel
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.72 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.885 2.065 2.115 2.065 2.115 2.58 3.28 2.58 3.51 2.58 3.51 2.12 4.4 2.12 4.4 2.35 3.77 2.35 3.77 2.81 3.28 2.81 1.885 2.81  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.81 2.12 1.435 2.12 1.435 3.04 3.28 3.04 4.43 3.04 4.43 2.89 4.66 2.89 4.66 2.12 5.47 2.12 5.47 2.35 4.89 2.35 4.89 3.27 3.28 3.27 1.205 3.27 1.205 2.35 0.81 2.35  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.675 3.5 5.305 3.5 5.305 2.58 5.75 2.58 5.75 1.37 4.69 1.37 4.69 1.14 6.01 1.14 6.01 2.81 5.535 2.81 5.535 3.73 3.905 3.73 3.905 4.31 3.675 4.31  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.285 4.59 0.285 3.5 0.515 3.5 0.515 4.59 2.325 4.59 2.325 3.5 2.555 3.5 2.555 4.59 3.28 4.59 5.765 4.59 5.765 3.5 5.995 3.5 5.995 4.59 6.15 4.59 6.72 4.59 6.72 5.49 6.15 5.49 3.28 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.72 -0.45 6.72 0.45 2.555 0.45 2.555 1.355 2.325 1.355 2.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.285 1.015 0.515 1.015 0.515 1.605 2.575 1.605 2.575 2.12 3.28 2.12 3.28 2.35 2.345 2.35 2.345 1.835 0.515 1.835 0.515 2.58 0.975 2.58 0.975 3.5 1.535 3.5 1.535 4.31 1.305 4.31 1.305 3.73 0.745 3.73 0.745 2.81 0.285 2.81  ;
        POLYGON 3.625 0.68 6.15 0.68 6.15 0.91 3.855 0.91 3.855 1.655 3.625 1.655  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.995 2 2.225 2 2.225 2.515 3.49 2.515 4.07 2.515 4.07 1.21 4.455 1.21 4.455 2.745 3.49 2.745 1.995 2.745  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.055 1.765 2.055 1.765 2.975 3.49 2.975 5.19 2.975 5.19 2.135 5.475 2.135 5.475 3.205 3.49 3.205 1.535 3.205 1.535 2.285 0.87 2.285  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 1.21 7.665 1.21 7.665 0.68 7.895 0.68 7.895 3.775 7.665 3.775 7.665 1.59 7.43 1.59  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.435 2.665 3.435 2.665 4.59 3.49 4.59 6.11 4.59 6.545 4.59 6.545 3.875 6.775 3.875 6.775 4.59 7.215 4.59 8.685 4.59 8.685 2.965 8.915 2.965 8.915 4.59 9.52 4.59 9.52 5.49 7.215 5.49 6.11 5.49 3.49 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 9.015 0.45 9.015 1.435 8.785 1.435 8.785 0.45 6.775 0.45 6.775 1.31 6.545 1.31 6.545 0.45 6.055 0.45 6.055 1.31 5.825 1.31 5.825 0.45 2.715 0.45 2.715 0.965 2.485 0.965 2.485 0.45 0.475 0.45 0.475 0.965 0.245 0.965 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.54 1.31 1.54 1.31 0.68 1.65 0.68 1.65 1.54 2.685 1.54 2.685 2.055 3.49 2.055 3.49 2.285 2.455 2.285 2.455 1.77 0.575 1.77 0.575 3.775 0.345 3.775  ;
        POLYGON 3.785 3.435 4.015 3.435 4.015 4.015 6.11 4.015 6.11 4.245 3.785 4.245  ;
        POLYGON 4.75 3.435 5.705 3.435 5.705 1.905 4.685 1.905 4.685 0.91 3.73 0.91 3.73 0.68 4.915 0.68 4.915 1.675 7.215 1.675 7.215 2.115 5.935 2.115 5.935 3.665 4.75 3.665  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.63 3.39 2.63 3.62 2.63 3.62 2.17 4.51 2.17 4.51 2.4 3.85 2.4 3.85 2.86 3.39 2.86 1.83 2.86  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.985 1.77 0.985 3.09 3.39 3.09 4.625 3.09 4.625 2.6 5.245 2.6 5.245 2.115 5.475 2.115 5.475 2.83 4.855 2.83 4.855 3.32 3.39 3.32 0.755 3.32 0.755 2.455 0.71 2.455  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 2.89 7.665 2.89 7.665 0.68 7.895 0.68 7.895 1.72 9.905 1.72 9.905 0.68 10.135 0.68 10.135 3.685 9.855 3.685 9.855 1.95 7.895 1.95 7.895 3.685 7.665 3.685 7.665 3.27 7.43 3.27  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.665 4.59 2.665 3.875 2.895 3.875 2.895 4.59 3.39 4.59 6.11 4.59 6.645 4.59 6.645 3.875 6.875 3.875 6.875 4.59 7.315 4.59 8.735 4.59 8.735 3.875 8.965 3.875 8.965 4.59 10.925 4.59 10.925 2.875 11.155 2.875 11.155 4.59 11.76 4.59 11.76 5.49 7.315 5.49 6.11 5.49 3.39 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 11.255 0.45 11.255 1.49 11.025 1.49 11.025 0.45 9.015 0.45 9.015 1.49 8.785 1.49 8.785 0.45 6.775 0.45 6.775 1.425 6.545 1.425 6.545 0.45 6.055 0.45 6.055 1.425 5.825 1.425 5.825 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 1.31 1.365 1.31 1.365 0.68 1.595 0.68 1.595 1.31 2.55 1.31 2.55 2.17 3.39 2.17 3.39 2.4 2.32 2.4 2.32 1.54 0.48 1.54 0.48 2.875 0.525 2.875 0.525 3.215 0.25 3.215  ;
        POLYGON 3.785 3.55 4.015 3.55 4.015 4.13 6.11 4.13 6.11 4.36 3.785 4.36  ;
        POLYGON 4.75 3.55 5.705 3.55 5.705 1.885 3.785 1.885 3.785 0.68 4.015 0.68 4.015 1.655 7.315 1.655 7.315 2.455 7.085 2.455 7.085 1.885 5.935 1.885 5.935 3.78 4.75 3.78  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.88 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.995 1.815 2.225 1.815 2.225 2.33 3.44 2.33 3.67 2.33 3.67 1.87 4.51 1.87 4.51 2.1 3.9 2.1 3.9 2.71 3.44 2.71 1.995 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 1.77 1.53 1.77 1.53 2.94 3.44 2.94 5.245 2.94 5.245 1.815 5.475 1.815 5.475 3.17 3.44 3.17 1.3 3.17 1.3 2.15 0.87 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.09 1.87 8.97 1.87 8.97 2.33 9.54 2.33 9.77 2.33 9.77 1.87 10.71 1.87 10.71 2.1 10 2.1 10 2.71 9.54 2.71 8.74 2.71 8.74 2.1 8.09 2.1  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9125 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.985 3.49 11.685 3.49 11.685 3.415 11.73 3.415 11.96 3.415 11.96 1.59 10.95 1.59 10.95 1.21 12.19 1.21 12.19 3.645 11.855 3.645 11.855 3.72 11.73 3.72 10.215 3.72 10.215 4.36 9.985 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.55 2.665 3.55 2.665 4.59 3.44 4.59 6.055 4.59 6.545 4.59 6.545 3.855 6.775 3.855 6.775 4.59 8.815 4.59 8.815 3.875 9.045 3.875 9.045 4.59 11.73 4.59 12.025 4.59 12.025 3.875 12.255 3.875 12.255 4.59 12.41 4.59 12.88 4.59 12.88 5.49 12.41 5.49 11.73 5.49 6.055 5.49 3.44 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.88 -0.45 12.88 0.45 8.815 0.45 8.815 1.08 8.585 1.08 8.585 0.45 6.055 0.45 6.055 1.08 5.825 1.08 5.825 0.45 2.715 0.45 2.715 1.08 2.485 1.08 2.485 0.45 0.475 0.45 0.475 1.08 0.245 1.08 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.31 1.365 1.31 1.365 0.74 1.595 0.74 1.595 1.31 2.685 1.31 2.685 1.87 3.44 1.87 3.44 2.1 2.455 2.1 2.455 1.54 0.575 1.54 0.575 3.89 0.345 3.89  ;
        POLYGON 3.785 3.55 4.015 3.55 4.015 4.13 5.825 4.13 5.825 3.855 6.055 3.855 6.055 4.36 3.785 4.36  ;
        POLYGON 6.545 1.04 6.775 1.04 6.775 1.41 9.54 1.41 9.54 2.1 9.2 2.1 9.2 1.64 7.795 1.64 7.795 3.64 7.565 3.64 7.565 1.64 6.545 1.64  ;
        POLYGON 5.955 3.395 7.235 3.395 7.235 3.87 8.355 3.87 8.355 3.03 11.285 3.03 11.285 1.87 11.73 1.87 11.73 2.1 11.515 2.1 11.515 3.26 8.585 3.26 8.585 4.1 7.005 4.1 7.005 3.625 5.775 3.625 5.775 3.63 5.035 3.63 5.035 3.89 4.805 3.89 4.805 3.4 5.725 3.4 5.725 1.54 3.785 1.54 3.785 0.74 4.015 0.74 4.015 1.31 5.955 1.31 5.955 1.87 7.27 1.87 7.27 2.1 5.955 2.1  ;
        POLYGON 9.885 0.74 12.41 0.74 12.41 0.97 10.115 0.97 10.115 1.55 9.885 1.55  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 1.72 4.33 1.72 4.33 2.18 4.575 2.18 4.575 2.52 4.07 2.52 4.07 1.95 2.395 1.95 2.395 2.52 2.165 2.52  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.025 2.18 1.255 2.18 1.255 3.21 3.555 3.21 5.19 3.21 5.19 2.18 5.595 2.18 5.595 3.44 3.555 3.44 1.025 3.44  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.31 2.77 9.86 2.77 10.23 2.77 10.23 2.31 10.93 2.31 10.93 2.54 10.49 2.54 10.49 3 9.86 3 8.31 3  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.772 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.015 3.155 13.685 3.155 13.915 3.155 13.915 1.945 12.965 1.945 12.965 0.845 13.29 0.845 13.29 1.715 15.205 1.715 15.205 0.845 15.435 0.845 15.435 1.945 14.145 1.945 14.145 3.155 15.385 3.155 15.385 4.36 15.155 4.36 15.155 3.385 13.685 3.385 13.245 3.385 13.245 4.36 13.015 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.605 4.59 2.605 3.67 2.835 3.67 2.835 4.59 3.555 4.59 6.23 4.59 8.805 4.59 8.805 3.615 9.035 3.615 9.035 4.59 9.86 4.59 12.475 4.59 13.685 4.59 14.035 4.59 14.035 3.615 14.265 3.615 14.265 4.59 15.68 4.59 15.68 5.49 13.685 5.49 12.475 5.49 9.86 5.49 6.23 5.49 3.555 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 14.315 0.45 14.315 1.485 14.085 1.485 14.085 0.45 12.475 0.45 12.475 1.16 12.245 1.16 12.245 0.45 9.315 0.45 9.315 1.18 9.085 1.18 9.085 0.45 6.895 0.45 6.895 1.185 6.665 1.185 6.665 0.45 6.175 0.45 6.175 1.185 5.945 1.185 5.945 0.45 2.835 0.45 2.835 1.185 2.605 1.185 2.605 0.45 0.595 0.45 0.595 1.185 0.365 1.185 0.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.465 1.72 1.485 1.72 1.485 0.845 1.715 0.845 1.715 2.75 3.325 2.75 3.325 2.18 3.555 2.18 3.555 2.98 1.485 2.98 1.485 1.95 0.695 1.95 0.695 3.955 0.465 3.955  ;
        POLYGON 3.905 3.67 4.135 3.67 4.135 4.13 6.23 4.13 6.23 4.36 3.905 4.36  ;
        POLYGON 6.765 2.75 7.785 2.75 7.785 1.145 8.015 1.145 8.015 2.31 9.86 2.31 9.86 2.54 8.015 2.54 8.015 2.98 6.995 2.98 6.995 4.36 6.765 4.36  ;
        POLYGON 4.87 3.67 5.825 3.67 5.825 2.29 7.205 2.29 7.205 1.645 4.55 1.645 4.55 1.13 3.85 1.13 3.85 0.9 4.78 0.9 4.78 1.415 7.205 1.415 7.205 0.685 8.475 0.685 8.475 1.85 11.895 1.85 11.895 2.52 11.665 2.52 11.665 2.08 8.245 2.08 8.245 0.915 7.435 0.915 7.435 2.52 6.055 2.52 6.055 3.9 4.87 3.9  ;
        POLYGON 10.15 3.55 12.475 3.55 12.475 4.36 12.245 4.36 12.245 3.9 10.15 3.9  ;
        POLYGON 11.17 2.93 12.125 2.93 12.125 1.62 10.205 1.62 10.205 0.845 10.435 0.845 10.435 1.39 12.355 1.39 12.355 2.18 13.685 2.18 13.685 2.52 12.355 2.52 12.355 3.16 11.17 3.16  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8595 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.99 1.77 4.33 1.77 4.33 2.395 3.99 2.395 3.99 2 2.33 2 2.33 2.36 1.99 2.36  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8595 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 2.11 1.19 2.11 1.19 3.05 3.29 3.05 3.51 3.05 3.51 2.89 3.74 2.89 3.74 2.625 5.01 2.625 5.01 2.165 5.35 2.165 5.35 2.855 3.97 2.855 3.97 3.28 3.29 3.28 0.96 3.28  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.145 2.775 9.785 2.775 10.23 2.775 10.23 2.33 10.805 2.33 10.805 2.56 10.49 2.56 10.49 3.005 9.785 3.005 8.145 3.005  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.593 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.94 3.415 13.665 3.415 13.895 3.415 13.895 2 12.84 2 12.84 0.845 13.07 0.845 13.07 1.77 15.08 1.77 15.08 0.845 15.31 0.845 15.31 1.885 17.32 1.885 17.32 0.845 17.55 0.845 17.55 4.345 17.22 4.345 17.22 2.115 15.26 2.115 15.26 4.345 15.03 4.345 15.03 2.15 14.125 2.15 14.125 3.645 13.665 3.645 13.17 3.645 13.17 4.345 12.94 4.345  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.535 2.615 3.535 2.615 4.59 3.29 4.59 6.11 4.59 8.64 4.59 8.64 3.535 8.87 3.535 8.87 4.59 9.785 4.59 12.35 4.59 13.665 4.59 13.96 4.59 13.96 3.875 14.19 3.875 14.19 4.59 16.15 4.59 16.15 3.875 16.38 3.875 16.38 4.59 17.92 4.59 17.92 5.49 13.665 5.49 12.35 5.49 9.785 5.49 6.11 5.49 3.29 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 16.43 0.45 16.43 1.655 16.2 1.655 16.2 0.45 14.19 0.45 14.19 1.165 13.96 1.165 13.96 0.45 12.35 0.45 12.35 1.165 12.12 1.165 12.12 0.45 9.19 0.45 9.19 1.165 8.96 1.165 8.96 0.45 5.645 0.45 5.645 0.845 6.73 0.845 6.73 1.48 6.5 1.48 6.5 1.185 5.415 1.185 5.415 0.45 2.715 0.45 2.715 1.185 2.485 1.185 2.485 0.45 0.475 0.45 0.475 1.185 0.245 1.185 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.65 1.365 1.65 1.365 0.845 1.65 0.845 1.65 2.59 3.29 2.59 3.29 2.82 1.42 2.82 1.42 1.88 0.575 1.88 0.575 3.875 0.345 3.875  ;
        POLYGON 3.605 3.535 3.835 3.535 3.835 4.105 5.88 4.105 5.88 3.535 6.11 3.535 6.11 4.335 3.605 4.335  ;
        POLYGON 6.6 2.68 7.62 2.68 7.62 1.14 7.85 1.14 7.85 2.315 9.785 2.315 9.785 2.545 7.85 2.545 7.85 2.91 6.83 2.91 6.83 3.875 6.6 3.875  ;
        POLYGON 4.625 3.085 5.58 3.085 5.58 1.935 4.56 1.935 4.56 1.13 3.55 1.13 3.55 0.9 4.79 0.9 4.79 1.705 5.63 1.705 5.63 1.71 7.04 1.71 7.04 0.68 8.31 0.68 8.31 1.855 11.825 1.855 11.825 2.085 8.08 2.085 8.08 0.91 7.27 0.91 7.27 2.45 7.04 2.45 7.04 1.94 5.81 1.94 5.81 3.315 4.855 3.315 4.855 3.875 4.625 3.875  ;
        POLYGON 10.08 3.55 10.31 3.55 10.31 4.13 12.12 4.13 12.12 3.55 12.35 3.55 12.35 4.36 10.08 4.36  ;
        POLYGON 11.1 2.315 12.055 2.315 12.055 1.625 10.08 1.625 10.08 0.815 10.31 0.815 10.31 1.395 12.285 1.395 12.285 2.23 13.665 2.23 13.665 2.545 11.33 2.545 11.33 3.9 11.1 3.9  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.72 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.905 2.87 1.905 2.87 2.33 3.44 2.33 3.885 2.33 3.885 1.85 4.455 1.85 4.455 2.19 4.115 2.19 4.115 2.71 3.44 2.71 2.64 2.71 2.64 2.135 1.94 2.135  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.85 1.015 1.85 1.015 2.94 3.44 2.94 4.345 2.94 4.345 2.47 4.83 2.47 4.83 1.905 5.53 1.905 5.53 2.135 5.06 2.135 5.06 2.7 4.575 2.7 4.575 3.17 3.44 3.17 0.71 3.17  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.805 3.04 5.19 3.04 5.19 2.89 5.76 2.89 5.76 1.62 3.785 1.62 3.785 0.81 4.015 0.81 4.015 1.39 5.99 1.39 5.99 3.12 5.45 3.12 5.45 3.27 5.035 3.27 5.035 3.9 4.805 3.9  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.4 2.665 3.4 2.665 4.59 3.44 4.59 6.055 4.59 6.72 4.59 6.72 5.49 6.055 5.49 3.44 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.72 -0.45 6.72 0.45 6.055 0.45 6.055 1.16 5.825 1.16 5.825 0.45 2.715 0.45 2.715 1.15 2.485 1.15 2.485 0.45 0.475 0.45 0.475 1.15 0.245 1.15 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 1.39 1.365 1.39 1.365 0.81 1.595 0.81 1.595 1.39 3.44 1.39 3.44 2.1 3.1 2.1 3.1 1.62 0.48 1.62 0.48 3.4 0.575 3.4 0.575 3.74 0.25 3.74  ;
        POLYGON 3.785 3.4 4.015 3.4 4.015 4.13 5.825 4.13 5.825 3.4 6.055 3.4 6.055 4.36 3.785 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 1.87 2.55 1.87 2.55 2.5 3.185 2.5 4.07 2.5 4.07 1.77 4.355 1.77 4.355 2.73 3.185 2.73 2.32 2.73 2.32 2.1 1.79 2.1  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.77 2.235 1.46 2.235 1.46 2.33 2.09 2.33 2.09 2.96 3.185 2.96 5.145 2.96 5.145 2.18 5.375 2.18 5.375 3.19 3.185 3.19 1.86 3.19 1.86 2.71 1.27 2.71 1.27 2.465 0.77 2.465  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 1.21 7.665 1.21 7.665 0.84 7.895 0.84 7.895 4.23 7.665 4.23 7.665 1.59 7.43 1.59  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.585 0.475 3.585 0.475 4.59 2.285 4.59 2.285 3.585 2.515 3.585 2.515 4.59 3.185 4.59 5.725 4.59 5.725 3.88 5.955 3.88 5.955 4.59 6.645 4.59 6.645 3.585 6.875 3.585 6.875 4.59 7.37 4.59 8.685 4.59 8.685 3.585 8.915 3.585 8.915 4.59 9.52 4.59 9.52 5.49 7.37 5.49 3.185 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 9.015 0.45 9.015 1.65 8.785 1.65 8.785 0.45 6.775 0.45 6.775 1.445 6.545 1.445 6.545 0.45 2.515 0.45 2.515 1.18 2.285 1.18 2.285 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.84 0.475 0.84 0.475 1.41 3.185 1.41 3.185 2.27 2.955 2.27 2.955 1.64 0.475 1.64 0.475 2.94 1.495 2.94 1.495 4.31 1.265 4.31 1.265 3.17 0.245 3.17  ;
        POLYGON 3.585 0.68 6.055 0.68 6.055 1.49 5.825 1.49 5.825 0.91 3.815 0.91 3.815 1.65 3.585 1.65  ;
        POLYGON 3.685 3.42 5.605 3.42 5.605 1.95 4.705 1.95 4.705 1.14 4.935 1.14 4.935 1.72 5.825 1.72 5.825 1.88 7.37 1.88 7.37 2.11 5.835 2.11 5.835 3.65 3.915 3.65 3.915 4.23 3.685 4.23  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 2.33 3.29 2.33 4.36 2.33 4.36 2.71 3.29 2.71 1.79 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.77 2.33 1.11 2.33 1.11 2.94 3.29 2.94 4.63 2.94 4.63 2.33 5.43 2.33 5.43 2.71 4.86 2.71 4.86 3.17 3.29 3.17 0.77 3.17  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 3.45 7.665 3.45 7.665 0.845 7.895 0.845 7.895 1.885 9.905 1.885 9.905 0.845 10.135 0.845 10.135 4.36 9.855 4.36 9.855 2.115 7.895 2.115 7.895 4.36 7.43 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.86 0.475 3.86 0.475 4.59 2.285 4.59 2.285 3.86 2.515 3.86 2.515 4.59 3.29 4.59 5.725 4.59 5.725 3.86 5.955 3.86 5.955 4.59 6.645 4.59 6.645 3.86 6.875 3.86 6.875 4.59 7.315 4.59 8.735 4.59 8.735 3.86 8.965 3.86 8.965 4.59 10.925 4.59 10.925 3.86 11.155 3.86 11.155 4.59 11.76 4.59 11.76 5.49 7.315 5.49 3.29 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 11.255 0.45 11.255 1.655 11.025 1.655 11.025 0.45 9.015 0.45 9.015 1.655 8.785 1.655 8.785 0.45 6.775 0.45 6.775 1.165 6.545 1.165 6.545 0.45 2.57 0.45 2.57 1.595 2.23 1.595 2.23 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 1.365 0.53 1.365 0.53 1.87 3.29 1.87 3.29 2.1 0.42 2.1 0.42 3.4 1.495 3.4 1.495 4.065 1.265 4.065 1.265 3.63 0.19 3.63  ;
        POLYGON 3.585 0.83 6.055 0.83 6.055 1.64 5.825 1.64 5.825 1.06 3.815 1.06 3.815 1.65 3.585 1.65  ;
        POLYGON 3.635 3.4 5.66 3.4 5.66 2.1 4.705 2.1 4.705 1.31 4.935 1.31 4.935 1.87 7.315 1.87 7.315 2.21 5.89 2.21 5.89 3.63 3.865 3.63 3.865 4.36 3.635 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_4
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.88 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.89 1.77 2.42 1.77 2.42 1.41 4.455 1.41 4.455 2.21 4.225 2.21 4.225 1.64 2.65 1.64 2.65 2.155 1.89 2.155  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.925 1.87 1.155 1.87 1.155 2.845 3.335 2.845 5.245 2.845 5.245 1.87 5.475 1.87 5.475 3.075 3.335 3.075 1.53 3.075 1.53 3.27 0.925 3.27  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.99 2.33 8.335 2.33 8.335 2.48 9.74 2.48 10.525 2.48 10.525 1.87 10.755 1.87 10.755 2.71 9.74 2.71 7.99 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.105 2.89 11.775 2.89 12.005 2.89 12.005 1.155 10.03 1.155 10.03 0.895 10.37 0.895 10.37 0.925 12.235 0.925 12.235 3.27 11.775 3.27 11.335 3.27 11.335 3.7 11.105 3.7  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.305 2.615 3.305 2.615 4.59 3.335 4.59 6.11 4.59 8.685 4.59 8.685 2.965 8.915 2.965 8.915 4.59 9.74 4.59 12.635 4.59 12.88 4.59 12.88 5.49 12.635 5.49 9.74 5.49 6.11 5.49 3.335 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.88 -0.45 12.88 0.45 12.355 0.45 12.355 0.695 12.125 0.695 12.125 0.45 9.015 0.45 9.015 1.18 8.785 1.18 8.785 0.45 6.775 0.45 6.775 1.18 6.545 1.18 6.545 0.45 6.055 0.45 6.055 1.18 5.825 1.18 5.825 0.45 2.715 0.45 2.715 1.18 2.485 1.18 2.485 0.45 0.475 0.45 0.475 1.18 0.245 1.18 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.41 1.365 1.41 1.365 0.84 1.615 0.84 1.615 2.385 3.105 2.385 3.105 1.87 3.335 1.87 3.335 2.615 1.385 2.615 1.385 1.64 0.575 1.64 0.575 3.645 0.345 3.645  ;
        POLYGON 3.785 3.305 4.015 3.305 4.015 3.83 6.11 3.83 6.11 4.115 3.785 4.115  ;
        POLYGON 6.63 2.44 7.53 2.44 7.53 1.89 7.665 1.89 7.665 1.14 7.895 1.14 7.895 1.87 9.74 1.87 9.74 2.155 9.4 2.155 9.4 2.1 7.76 2.1 7.76 2.67 6.86 2.67 6.86 3.775 6.63 3.775  ;
        POLYGON 4.75 3.36 5.705 3.36 5.705 1.64 4.685 1.64 4.685 1.125 3.73 1.125 3.73 0.895 4.915 0.895 4.915 1.41 7.205 1.41 7.205 0.68 8.555 0.68 8.555 1.41 11.775 1.41 11.775 2.21 11.545 2.21 11.545 1.64 8.325 1.64 8.325 0.91 7.435 0.91 7.435 1.62 7.3 1.62 7.3 2.21 7.07 2.21 7.07 1.64 5.935 1.64 5.935 3.59 4.75 3.59  ;
        POLYGON 10.085 3.305 10.315 3.305 10.315 4.005 12.405 4.005 12.405 3.425 12.635 3.425 12.635 4.235 10.085 4.235  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_1
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.51 4.455 1.51 4.455 2.025 4.225 2.025 4.225 1.74 2.17 1.74 2.17 2.2 1.83 2.2  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.91 1.915 1.14 1.915 1.14 2.89 3.44 2.89 3.67 2.89 3.67 2.255 5.19 2.255 5.19 1.97 5.53 1.97 5.53 2.485 3.9 2.485 3.9 3.27 3.44 3.27 0.91 3.27  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.09 2.37 9.54 2.37 9.67 2.37 9.67 2.33 10.71 2.33 10.71 2.71 9.54 2.71 8.09 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.772 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.845 3.415 13.57 3.415 13.8 3.415 13.8 1.67 12.845 1.67 12.845 0.845 13.29 0.845 13.29 1.44 15.085 1.44 15.085 0.845 15.315 0.845 15.315 3.685 14.985 3.685 14.985 1.67 14.03 1.67 14.03 3.645 13.57 3.645 13.075 3.645 13.075 4.32 12.845 4.32  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.51 2.665 3.51 2.665 4.59 3.44 4.59 6.055 4.59 6.545 4.59 6.545 3.45 6.775 3.45 6.775 4.59 8.815 4.59 8.815 4.35 9.045 4.35 9.045 4.59 12.025 4.59 12.025 4.35 12.255 4.35 12.255 4.59 13.57 4.59 13.865 4.59 13.865 3.875 14.095 3.875 14.095 4.59 15.68 4.59 15.68 5.49 13.57 5.49 6.055 5.49 3.44 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 14.195 0.45 14.195 1.165 13.965 1.165 13.965 0.45 8.815 0.45 8.815 1.185 8.585 1.185 8.585 0.45 6.055 0.45 6.055 1.185 5.825 1.185 5.825 0.45 2.715 0.45 2.715 1.185 2.485 1.185 2.485 0.45 0.475 0.45 0.475 1.185 0.245 1.185 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.455 1.365 1.455 1.365 0.845 1.6 0.845 1.6 2.43 3.1 2.43 3.1 1.97 3.44 1.97 3.44 2.66 1.37 2.66 1.37 1.685 0.575 1.685 0.575 3.85 0.345 3.85  ;
        POLYGON 3.785 3.51 4.015 3.51 4.015 4.13 5.825 4.13 5.825 3.175 6.055 3.175 6.055 4.36 3.785 4.36  ;
        POLYGON 6.49 0.9 7.795 0.9 7.795 1.91 9.54 1.91 9.54 2.14 7.795 2.14 7.795 3.235 7.565 3.235 7.565 1.13 6.49 1.13  ;
        POLYGON 4.805 2.715 7.005 2.715 7.005 1.645 4.685 1.645 4.685 1.13 3.73 1.13 3.73 0.9 4.915 0.9 4.915 1.415 7.235 1.415 7.235 3.465 10.94 3.465 10.94 2.18 11.73 2.18 11.73 2.41 11.17 2.41 11.17 3.695 7.005 3.695 7.005 2.945 5.035 2.945 5.035 3.9 4.805 3.9  ;
        POLYGON 9.885 0.68 12.355 0.68 12.355 1.49 12.125 1.49 12.125 0.91 10.115 0.91 10.115 1.655 9.885 1.655  ;
        POLYGON 9.93 3.925 11.265 3.925 11.265 3.905 11.71 3.905 11.71 2.64 11.96 2.64 11.96 1.95 11.005 1.95 11.005 1.14 11.235 1.14 11.235 1.72 12.185 1.72 12.185 1.9 13.57 1.9 13.57 2.13 12.19 2.13 12.19 2.87 11.94 2.87 11.94 4.135 11.36 4.135 11.36 4.155 9.93 4.155  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_2
#--------EOF---------

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8595 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.21 2.09 1.21 2.09 1.775 4.275 1.775 4.275 2.52 4.045 2.52 4.045 2.005 2.17 2.005 2.17 2.135 1.83 2.135  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8595 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.905 2.18 1.135 2.18 1.135 2.825 2.735 2.825 2.735 2.775 3.31 2.775 4.63 2.775 4.63 2.18 5.295 2.18 5.295 2.71 4.86 2.71 4.86 3.005 3.31 3.005 2.88 3.005 2.88 3.055 0.905 3.055  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.91 2.475 9.41 2.475 9.67 2.475 9.67 2.33 10.48 2.33 10.48 2.71 9.41 2.71 7.91 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.593 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.765 3.235 13.49 3.235 13.72 3.235 13.72 1.72 13.59 1.72 13.59 1.49 12.665 1.49 12.665 0.68 12.895 0.68 12.895 1.21 14.905 1.21 14.905 0.845 15.135 0.845 15.135 1.885 17.145 1.885 17.145 0.845 17.375 0.845 17.375 4.36 17.045 4.36 17.045 2.115 15.185 2.115 15.185 4.36 14.955 4.36 14.955 2.03 13.95 2.03 13.95 3.465 13.49 3.465 12.995 3.465 12.995 4.36 12.765 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.695 2.615 3.695 2.615 4.59 3.31 4.59 5.875 4.59 6.365 4.59 6.365 3.015 6.595 3.015 6.595 4.59 8.685 4.59 8.685 3.865 8.915 3.865 8.915 4.59 11.845 4.59 11.845 4.35 12.075 4.35 12.075 4.59 13.49 4.59 13.785 4.59 13.785 3.695 14.015 3.695 14.015 4.59 15.975 4.59 15.975 3.695 16.205 3.695 16.205 4.59 17.92 4.59 17.92 5.49 13.49 5.49 5.875 5.49 3.31 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 16.255 0.45 16.255 1.655 16.025 1.655 16.025 0.45 14.015 0.45 14.015 0.695 13.785 0.695 13.785 0.45 8.635 0.45 8.635 1.185 8.405 1.185 8.405 0.45 5.875 0.45 5.875 1.185 5.645 1.185 5.645 0.45 2.715 0.45 2.715 1.185 2.485 1.185 2.485 0.45 0.475 0.45 0.475 1.185 0.245 1.185 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.72 1.365 1.72 1.365 0.845 1.595 0.845 1.595 2.365 2.38 2.365 2.38 2.235 3.31 2.235 3.31 2.465 2.59 2.465 2.59 2.595 1.365 2.595 1.365 1.95 0.575 1.95 0.575 4.035 0.345 4.035  ;
        POLYGON 3.605 3.695 3.835 3.695 3.835 4.13 5.645 4.13 5.645 3.695 5.875 3.695 5.875 4.36 3.605 4.36  ;
        POLYGON 6.365 0.845 6.595 0.845 6.595 1.72 7.615 1.72 7.615 2.015 9.41 2.015 9.41 2.245 7.615 2.245 7.615 3.22 7.385 3.22 7.385 1.95 6.365 1.95  ;
        POLYGON 4.625 3.235 5.525 3.235 5.525 1.645 4.465 1.645 4.465 1.13 3.55 1.13 3.55 0.9 4.695 0.9 4.695 1.415 5.755 1.415 5.755 2.18 7.055 2.18 7.055 3.45 8.405 3.45 8.405 3.405 11.265 3.405 11.265 2.18 11.495 2.18 11.495 3.635 8.545 3.635 8.545 3.68 6.825 3.68 6.825 2.41 5.755 2.41 5.755 3.465 4.855 3.465 4.855 3.9 4.625 3.9  ;
        POLYGON 9.705 0.68 12.175 0.68 12.175 1.49 11.945 1.49 11.945 0.91 9.935 0.91 9.935 1.655 9.705 1.655  ;
        POLYGON 9.7 3.865 11.725 3.865 11.725 1.95 10.825 1.95 10.825 1.315 11.055 1.315 11.055 1.72 11.955 1.72 11.955 1.93 13.49 1.93 13.49 2.16 11.955 2.16 11.955 4.095 9.7 4.095  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_4
#--------EOF---------


END LIBRARY
