magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 4902 1094
<< pwell >>
rect -86 -86 4902 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
rect 1468 69 1588 333
rect 1692 69 1812 333
rect 2060 69 2180 333
rect 2284 69 2404 333
rect 2508 69 2628 333
rect 2732 69 2852 333
rect 2956 69 3076 333
rect 3180 69 3300 333
rect 3404 69 3524 333
rect 3628 69 3748 333
rect 3852 69 3972 333
rect 4076 69 4196 333
rect 4300 69 4420 333
rect 4524 69 4644 333
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 806 573 906 939
rect 1030 573 1130 939
rect 1254 573 1354 939
rect 1478 573 1578 939
rect 1702 573 1802 939
rect 2060 647 2160 939
rect 2304 647 2404 939
rect 2508 647 2608 939
rect 2732 647 2832 939
rect 2976 573 3076 939
rect 3190 573 3290 939
rect 3424 573 3524 939
rect 3638 573 3738 939
rect 3862 573 3962 939
rect 4086 573 4186 939
rect 4310 573 4410 939
rect 4524 573 4624 939
<< mvndiff >>
rect 36 291 124 333
rect 36 151 49 291
rect 95 151 124 291
rect 36 69 124 151
rect 244 291 348 333
rect 244 151 273 291
rect 319 151 348 291
rect 244 69 348 151
rect 468 291 572 333
rect 468 151 497 291
rect 543 151 572 291
rect 468 69 572 151
rect 692 291 796 333
rect 692 151 721 291
rect 767 151 796 291
rect 692 69 796 151
rect 916 197 1020 333
rect 916 151 945 197
rect 991 151 1020 197
rect 916 69 1020 151
rect 1140 291 1244 333
rect 1140 151 1169 291
rect 1215 151 1244 291
rect 1140 69 1244 151
rect 1364 197 1468 333
rect 1364 151 1393 197
rect 1439 151 1468 197
rect 1364 69 1468 151
rect 1588 291 1692 333
rect 1588 151 1617 291
rect 1663 151 1692 291
rect 1588 69 1692 151
rect 1812 197 1900 333
rect 1812 151 1841 197
rect 1887 151 1900 197
rect 1812 69 1900 151
rect 1972 197 2060 333
rect 1972 151 1985 197
rect 2031 151 2060 197
rect 1972 69 2060 151
rect 2180 274 2284 333
rect 2180 228 2209 274
rect 2255 228 2284 274
rect 2180 69 2284 228
rect 2404 197 2508 333
rect 2404 151 2433 197
rect 2479 151 2508 197
rect 2404 69 2508 151
rect 2628 285 2732 333
rect 2628 239 2657 285
rect 2703 239 2732 285
rect 2628 69 2732 239
rect 2852 197 2956 333
rect 2852 151 2881 197
rect 2927 151 2956 197
rect 2852 69 2956 151
rect 3076 285 3180 333
rect 3076 239 3105 285
rect 3151 239 3180 285
rect 3076 69 3180 239
rect 3300 197 3404 333
rect 3300 151 3329 197
rect 3375 151 3404 197
rect 3300 69 3404 151
rect 3524 274 3628 333
rect 3524 228 3553 274
rect 3599 228 3628 274
rect 3524 69 3628 228
rect 3748 197 3852 333
rect 3748 151 3777 197
rect 3823 151 3852 197
rect 3748 69 3852 151
rect 3972 285 4076 333
rect 3972 239 4001 285
rect 4047 239 4076 285
rect 3972 69 4076 239
rect 4196 291 4300 333
rect 4196 151 4225 291
rect 4271 151 4300 291
rect 4196 69 4300 151
rect 4420 285 4524 333
rect 4420 239 4449 285
rect 4495 239 4524 285
rect 4420 69 4524 239
rect 4644 291 4732 333
rect 4644 151 4673 291
rect 4719 151 4732 291
rect 4644 69 4732 151
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 358 939
rect 458 881 582 939
rect 458 741 487 881
rect 533 741 582 881
rect 458 573 582 741
rect 682 573 806 939
rect 906 861 1030 939
rect 906 721 935 861
rect 981 721 1030 861
rect 906 573 1030 721
rect 1130 573 1254 939
rect 1354 849 1478 939
rect 1354 803 1383 849
rect 1429 803 1478 849
rect 1354 573 1478 803
rect 1578 573 1702 939
rect 1802 861 2060 939
rect 1802 721 1831 861
rect 1877 721 2060 861
rect 1802 647 2060 721
rect 2160 849 2304 939
rect 2160 803 2189 849
rect 2235 803 2304 849
rect 2160 647 2304 803
rect 2404 861 2508 939
rect 2404 721 2433 861
rect 2479 721 2508 861
rect 2404 647 2508 721
rect 2608 849 2732 939
rect 2608 803 2637 849
rect 2683 803 2732 849
rect 2608 647 2732 803
rect 2832 861 2976 939
rect 2832 721 2861 861
rect 2907 721 2976 861
rect 2832 647 2976 721
rect 1802 573 1882 647
rect 2896 573 2976 647
rect 3076 573 3190 939
rect 3290 849 3424 939
rect 3290 803 3319 849
rect 3365 803 3424 849
rect 3290 573 3424 803
rect 3524 573 3638 939
rect 3738 861 3862 939
rect 3738 721 3767 861
rect 3813 721 3862 861
rect 3738 573 3862 721
rect 3962 573 4086 939
rect 4186 849 4310 939
rect 4186 803 4215 849
rect 4261 803 4310 849
rect 4186 573 4310 803
rect 4410 573 4524 939
rect 4624 861 4712 939
rect 4624 721 4653 861
rect 4699 721 4712 861
rect 4624 573 4712 721
<< mvndiffc >>
rect 49 151 95 291
rect 273 151 319 291
rect 497 151 543 291
rect 721 151 767 291
rect 945 151 991 197
rect 1169 151 1215 291
rect 1393 151 1439 197
rect 1617 151 1663 291
rect 1841 151 1887 197
rect 1985 151 2031 197
rect 2209 228 2255 274
rect 2433 151 2479 197
rect 2657 239 2703 285
rect 2881 151 2927 197
rect 3105 239 3151 285
rect 3329 151 3375 197
rect 3553 228 3599 274
rect 3777 151 3823 197
rect 4001 239 4047 285
rect 4225 151 4271 291
rect 4449 239 4495 285
rect 4673 151 4719 291
<< mvpdiffc >>
rect 69 721 115 861
rect 487 741 533 881
rect 935 721 981 861
rect 1383 803 1429 849
rect 1831 721 1877 861
rect 2189 803 2235 849
rect 2433 721 2479 861
rect 2637 803 2683 849
rect 2861 721 2907 861
rect 3319 803 3365 849
rect 3767 721 3813 861
rect 4215 803 4261 849
rect 4653 721 4699 861
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 806 939 906 983
rect 1030 939 1130 983
rect 1254 939 1354 983
rect 1478 939 1578 983
rect 1702 939 1802 983
rect 2060 939 2160 983
rect 2304 939 2404 983
rect 2508 939 2608 983
rect 2732 939 2832 983
rect 2976 939 3076 983
rect 3190 939 3290 983
rect 3424 939 3524 983
rect 3638 939 3738 983
rect 3862 939 3962 983
rect 4086 939 4186 983
rect 4310 939 4410 983
rect 4524 939 4624 983
rect 144 500 244 573
rect 144 454 185 500
rect 231 454 244 500
rect 144 377 244 454
rect 358 513 458 573
rect 582 513 682 573
rect 358 500 682 513
rect 358 454 623 500
rect 669 454 682 500
rect 358 441 682 454
rect 358 377 468 441
rect 124 333 244 377
rect 348 333 468 377
rect 572 377 682 441
rect 806 513 906 573
rect 1030 513 1130 573
rect 806 500 1130 513
rect 806 454 825 500
rect 871 454 1130 500
rect 806 441 1130 454
rect 806 377 916 441
rect 572 333 692 377
rect 796 333 916 377
rect 1020 377 1130 441
rect 1254 513 1354 573
rect 1478 513 1578 573
rect 1254 500 1578 513
rect 1254 454 1267 500
rect 1313 454 1578 500
rect 1254 441 1578 454
rect 1254 377 1364 441
rect 1020 333 1140 377
rect 1244 333 1364 377
rect 1468 377 1578 441
rect 1702 500 1802 573
rect 1702 454 1715 500
rect 1761 454 1802 500
rect 1702 377 1802 454
rect 2060 513 2160 647
rect 2304 513 2404 647
rect 2508 513 2608 647
rect 2732 513 2832 647
rect 2060 500 2832 513
rect 2060 454 2209 500
rect 2255 454 2433 500
rect 2479 454 2657 500
rect 2703 454 2832 500
rect 2060 441 2832 454
rect 1468 333 1588 377
rect 1692 333 1812 377
rect 2060 333 2180 441
rect 2284 333 2404 441
rect 2508 333 2628 441
rect 2732 377 2832 441
rect 2976 500 3076 573
rect 2976 454 3017 500
rect 3063 454 3076 500
rect 2976 377 3076 454
rect 3190 513 3290 573
rect 3424 513 3524 573
rect 3190 500 3524 513
rect 3190 454 3465 500
rect 3511 454 3524 500
rect 3190 441 3524 454
rect 3190 377 3300 441
rect 2732 333 2852 377
rect 2956 333 3076 377
rect 3180 333 3300 377
rect 3404 333 3524 441
rect 3638 513 3738 573
rect 3862 513 3962 573
rect 4086 513 4186 573
rect 4310 513 4410 573
rect 3638 500 3962 513
rect 3638 454 3828 500
rect 3874 454 3962 500
rect 3638 441 3962 454
rect 3638 377 3748 441
rect 3628 333 3748 377
rect 3852 377 3962 441
rect 4076 500 4410 513
rect 4076 454 4089 500
rect 4135 454 4410 500
rect 4076 441 4410 454
rect 3852 333 3972 377
rect 4076 333 4196 441
rect 4300 377 4410 441
rect 4524 500 4624 573
rect 4524 454 4537 500
rect 4583 454 4624 500
rect 4524 377 4624 454
rect 4300 333 4420 377
rect 4524 333 4644 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1468 25 1588 69
rect 1692 25 1812 69
rect 2060 25 2180 69
rect 2284 25 2404 69
rect 2508 25 2628 69
rect 2732 25 2852 69
rect 2956 25 3076 69
rect 3180 25 3300 69
rect 3404 25 3524 69
rect 3628 25 3748 69
rect 3852 25 3972 69
rect 4076 25 4196 69
rect 4300 25 4420 69
rect 4524 25 4644 69
<< polycontact >>
rect 185 454 231 500
rect 623 454 669 500
rect 825 454 871 500
rect 1267 454 1313 500
rect 1715 454 1761 500
rect 2209 454 2255 500
rect 2433 454 2479 500
rect 2657 454 2703 500
rect 3017 454 3063 500
rect 3465 454 3511 500
rect 3828 454 3874 500
rect 4089 454 4135 500
rect 4537 454 4583 500
<< metal1 >>
rect 0 918 4816 1098
rect 487 881 533 918
rect 69 861 115 872
rect 487 730 533 741
rect 935 861 981 872
rect 69 684 115 721
rect 1383 849 1429 918
rect 1383 792 1429 803
rect 1831 861 1877 872
rect 981 721 1831 746
rect 2189 849 2235 918
rect 2189 792 2235 803
rect 2433 861 2479 872
rect 1877 721 2433 746
rect 2637 849 2683 918
rect 2637 792 2683 803
rect 2861 861 2907 872
rect 2479 721 2861 746
rect 3319 849 3365 918
rect 3319 792 3365 803
rect 3714 861 3813 872
rect 3714 746 3767 861
rect 2907 721 3767 746
rect 4215 849 4261 918
rect 4215 792 4261 803
rect 4653 861 4699 872
rect 3813 721 4653 746
rect 935 700 4699 721
rect 935 684 981 700
rect 69 638 981 684
rect 3006 608 4238 654
rect 174 546 1416 592
rect 174 500 242 546
rect 814 500 882 546
rect 1370 500 1416 546
rect 2198 500 2714 542
rect 174 454 185 500
rect 231 454 242 500
rect 612 454 623 500
rect 669 454 726 500
rect 814 454 825 500
rect 871 454 882 500
rect 928 454 1267 500
rect 1313 454 1324 500
rect 1370 454 1715 500
rect 1761 454 1772 500
rect 2198 454 2209 500
rect 2255 454 2433 500
rect 2479 454 2657 500
rect 2703 454 2714 500
rect 3006 500 3074 608
rect 3828 578 4238 608
rect 3828 500 3874 578
rect 4192 500 4238 578
rect 3006 454 3017 500
rect 3063 454 3074 500
rect 3454 454 3465 500
rect 3511 454 3554 500
rect 680 435 726 454
rect 680 408 772 435
rect 928 408 974 454
rect 680 404 974 408
rect 273 348 635 394
rect 692 354 974 404
rect 3502 397 3554 454
rect 3828 443 3874 454
rect 3920 454 4089 500
rect 4135 454 4146 500
rect 4192 454 4537 500
rect 4583 454 4594 500
rect 3920 397 3966 454
rect 3502 351 3966 397
rect 4640 394 4699 700
rect 49 291 95 302
rect 49 90 95 151
rect 273 291 319 348
rect 589 302 635 348
rect 4012 348 4699 394
rect 4012 304 4058 348
rect 273 140 319 151
rect 497 291 543 302
rect 589 291 2703 302
rect 589 256 721 291
rect 497 90 543 151
rect 767 256 1169 291
rect 721 140 767 151
rect 945 197 991 208
rect 945 90 991 151
rect 1215 256 1617 291
rect 1169 140 1215 151
rect 1393 197 1439 208
rect 1393 90 1439 151
rect 1663 285 2703 291
rect 1663 274 2657 285
rect 1663 256 2209 274
rect 2198 228 2209 256
rect 2255 256 2657 274
rect 2255 228 2266 256
rect 2657 228 2703 239
rect 3105 285 4058 304
rect 3151 274 4001 285
rect 3151 258 3553 274
rect 3105 228 3151 239
rect 3542 228 3553 258
rect 3599 258 4001 274
rect 3599 228 3610 258
rect 4047 239 4058 285
rect 4001 228 4058 239
rect 4225 291 4271 302
rect 1617 140 1663 151
rect 1841 197 1887 208
rect 1841 90 1887 151
rect 1985 197 2031 208
rect 2422 182 2433 197
rect 2031 151 2433 182
rect 2479 182 2490 197
rect 2870 182 2881 197
rect 2479 151 2881 182
rect 2927 182 2938 197
rect 3318 182 3329 197
rect 2927 151 3329 182
rect 3375 182 3386 197
rect 3766 182 3777 197
rect 3375 151 3777 182
rect 3823 182 3834 197
rect 3823 151 4225 182
rect 4449 285 4495 348
rect 4449 228 4495 239
rect 4673 291 4719 302
rect 4271 151 4673 182
rect 1985 136 4719 151
rect 0 -90 4816 90
<< labels >>
flabel metal1 s 3006 608 4238 654 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 3920 454 4146 500 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 174 546 1416 592 0 FreeSans 200 0 0 0 B1
port 3 nsew default input
flabel metal1 s 928 454 1324 500 0 FreeSans 200 0 0 0 B2
port 4 nsew default input
flabel metal1 s 2198 454 2714 542 0 FreeSans 200 0 0 0 C
port 5 nsew default input
flabel metal1 s 0 918 4816 1098 0 FreeSans 200 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 497 208 543 302 0 FreeSans 200 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel metal1 s 4653 746 4699 872 0 FreeSans 200 0 0 0 ZN
port 6 nsew default output
rlabel metal1 s 3828 578 4238 608 1 A1
port 1 nsew default input
rlabel metal1 s 3006 578 3074 608 1 A1
port 1 nsew default input
rlabel metal1 s 4192 500 4238 578 1 A1
port 1 nsew default input
rlabel metal1 s 3828 500 3874 578 1 A1
port 1 nsew default input
rlabel metal1 s 3006 500 3074 578 1 A1
port 1 nsew default input
rlabel metal1 s 4192 454 4594 500 1 A1
port 1 nsew default input
rlabel metal1 s 3828 454 3874 500 1 A1
port 1 nsew default input
rlabel metal1 s 3006 454 3074 500 1 A1
port 1 nsew default input
rlabel metal1 s 3828 443 3874 454 1 A1
port 1 nsew default input
rlabel metal1 s 3454 454 3554 500 1 A2
port 2 nsew default input
rlabel metal1 s 3920 397 3966 454 1 A2
port 2 nsew default input
rlabel metal1 s 3502 397 3554 454 1 A2
port 2 nsew default input
rlabel metal1 s 3502 351 3966 397 1 A2
port 2 nsew default input
rlabel metal1 s 1370 500 1416 546 1 B1
port 3 nsew default input
rlabel metal1 s 814 500 882 546 1 B1
port 3 nsew default input
rlabel metal1 s 174 500 242 546 1 B1
port 3 nsew default input
rlabel metal1 s 1370 454 1772 500 1 B1
port 3 nsew default input
rlabel metal1 s 814 454 882 500 1 B1
port 3 nsew default input
rlabel metal1 s 174 454 242 500 1 B1
port 3 nsew default input
rlabel metal1 s 612 454 726 500 1 B2
port 4 nsew default input
rlabel metal1 s 928 435 974 454 1 B2
port 4 nsew default input
rlabel metal1 s 680 435 726 454 1 B2
port 4 nsew default input
rlabel metal1 s 928 408 974 435 1 B2
port 4 nsew default input
rlabel metal1 s 680 408 772 435 1 B2
port 4 nsew default input
rlabel metal1 s 680 404 974 408 1 B2
port 4 nsew default input
rlabel metal1 s 692 354 974 404 1 B2
port 4 nsew default input
rlabel metal1 s 3714 746 3813 872 1 ZN
port 6 nsew default output
rlabel metal1 s 2861 746 2907 872 1 ZN
port 6 nsew default output
rlabel metal1 s 2433 746 2479 872 1 ZN
port 6 nsew default output
rlabel metal1 s 1831 746 1877 872 1 ZN
port 6 nsew default output
rlabel metal1 s 935 746 981 872 1 ZN
port 6 nsew default output
rlabel metal1 s 69 746 115 872 1 ZN
port 6 nsew default output
rlabel metal1 s 935 700 4699 746 1 ZN
port 6 nsew default output
rlabel metal1 s 69 700 115 746 1 ZN
port 6 nsew default output
rlabel metal1 s 4640 684 4699 700 1 ZN
port 6 nsew default output
rlabel metal1 s 935 684 981 700 1 ZN
port 6 nsew default output
rlabel metal1 s 69 684 115 700 1 ZN
port 6 nsew default output
rlabel metal1 s 4640 638 4699 684 1 ZN
port 6 nsew default output
rlabel metal1 s 69 638 981 684 1 ZN
port 6 nsew default output
rlabel metal1 s 4640 394 4699 638 1 ZN
port 6 nsew default output
rlabel metal1 s 4012 348 4699 394 1 ZN
port 6 nsew default output
rlabel metal1 s 4449 304 4495 348 1 ZN
port 6 nsew default output
rlabel metal1 s 4012 304 4058 348 1 ZN
port 6 nsew default output
rlabel metal1 s 4449 258 4495 304 1 ZN
port 6 nsew default output
rlabel metal1 s 3105 258 4058 304 1 ZN
port 6 nsew default output
rlabel metal1 s 4449 228 4495 258 1 ZN
port 6 nsew default output
rlabel metal1 s 4001 228 4058 258 1 ZN
port 6 nsew default output
rlabel metal1 s 3542 228 3610 258 1 ZN
port 6 nsew default output
rlabel metal1 s 3105 228 3151 258 1 ZN
port 6 nsew default output
rlabel metal1 s 4215 792 4261 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3319 792 3365 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2637 792 2683 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2189 792 2235 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1383 792 1429 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 487 792 533 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 487 730 533 792 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 49 208 95 302 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1841 90 1887 208 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 208 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 208 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 208 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 208 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4816 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4816 1008
string GDS_END 234902
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 225688
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
