// This is the unpowered netlist.
module ffra (clk,
    rst,
    a,
    b,
    ci,
    o);
 input clk;
 input rst;
 input [7:0] a;
 input [7:0] b;
 input [15:0] ci;
 output [15:0] o;

 wire net2;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net1;

 gf180mcu_osu_sc_gp9t3v3__tiel ffra_2 (.Y(net2));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_3 (.Y(net3));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_4 (.Y(net4));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_5 (.Y(net5));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_6 (.Y(net6));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_7 (.Y(net7));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_8 (.Y(net8));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_9 (.Y(net9));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_10 (.Y(net10));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_11 (.Y(net11));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_12 (.Y(net12));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_13 (.Y(net13));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_14 (.Y(net14));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_15 (.Y(net15));
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_16 (.Y(net16));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_0 ();
 gf180mcu_osu_sc_gp9t3v3__tiel ffra_1 (.Y(net1));
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_0_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_1_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_2_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_3_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_4_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_5_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_6_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_7_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_8_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_9_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_10_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_11_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_12_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_13_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_14_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_15_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_16_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_17_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_18_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_19_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_20_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_21_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_22_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_23_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_24_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_25_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_26_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_27_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_28_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_29_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_30_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_31_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_32_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_33_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_34_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_35_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_36_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_37_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_38_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_39_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_40_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_41_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_42_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_43_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_44_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_45_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_46_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_47_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_48_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_49_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_50_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_51_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_52_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_53_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_54_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_55_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_56_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_57_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_58_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_59_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_60_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_61_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_62_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_63_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_64_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_65_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_66_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_67_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_68_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_69_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_70_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_71_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_72_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_73_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_74_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_75_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_76_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_77_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_78_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_79_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_80_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_81_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_82_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_83_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_84_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_85_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_86_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_1984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_2992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_3984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_4992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_5984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6976 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_6992 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7008 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7024 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7040 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7056 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7072 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7088 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7104 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7120 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7136 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7152 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7168 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7184 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7200 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7216 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7232 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7248 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7264 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7280 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7296 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7312 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7328 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7344 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7360 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7376 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7392 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7408 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7424 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7440 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7456 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7472 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7488 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7504 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7520 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7536 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7552 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7568 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7584 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7600 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7616 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7632 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7648 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7664 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7680 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7696 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7712 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7728 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7744 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7760 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7776 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7792 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7808 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7824 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7840 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7856 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7872 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7888 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7904 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7920 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7936 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7952 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7968 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_7984 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8000 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8016 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8032 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8048 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8064 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8080 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8096 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8288 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8304 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8320 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8336 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8352 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8368 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8384 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8400 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8416 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8432 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8448 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8464 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8480 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8496 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8512 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8528 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8544 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8560 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8576 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8592 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8608 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8624 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8640 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8656 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8672 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8688 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8704 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8720 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8736 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8752 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8768 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8784 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8800 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8816 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8832 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8848 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8864 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8880 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8896 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8912 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8928 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8944 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_87_8960 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_0 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_16 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_32 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_48 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_64 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_80 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_96 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_112 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_128 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_144 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_160 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_176 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_192 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_208 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_224 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_240 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_256 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_272 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_310 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_326 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_342 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_358 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_374 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_390 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_406 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_422 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_438 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_454 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_470 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_486 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_502 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_518 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_534 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_550 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_566 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_582 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_598 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_614 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_630 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_646 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_662 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_678 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_694 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_710 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_726 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_742 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_758 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_774 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_790 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_806 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_822 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_838 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_846 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_870 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_886 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_902 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_918 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_934 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_950 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_966 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_982 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_998 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1014 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1030 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1046 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1062 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1078 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1094 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1110 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1126 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1142 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1158 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1174 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1190 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1206 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1222 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1238 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1254 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1270 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1286 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1302 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1318 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1334 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1350 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1366 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1382 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_1398 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_1406 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1430 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1446 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1462 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1478 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1494 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1510 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1526 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1542 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1558 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1574 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1590 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1606 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1622 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1638 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1654 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1670 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1686 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1702 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1718 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1734 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1750 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1766 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1782 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1798 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1814 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1830 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1846 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1862 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1878 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1894 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1910 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1926 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1942 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_1958 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_1966 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_1990 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2006 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2022 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2038 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2054 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2070 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2086 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2102 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2118 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2134 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2150 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2166 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2182 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2198 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2214 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2230 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2246 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2262 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2278 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2294 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2310 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2326 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2342 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2358 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2374 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2390 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2406 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2422 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2438 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2454 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2470 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2486 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2502 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_2518 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_2526 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2550 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2566 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2582 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2598 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2614 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2630 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2646 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2662 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2678 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2694 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2710 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2726 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2742 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2758 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2774 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2790 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2806 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2822 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2838 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2854 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2870 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2886 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2902 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2918 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2934 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2950 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2966 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2982 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_2998 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3014 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3030 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3046 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3062 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_3078 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_3086 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3110 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3126 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3142 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3158 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3174 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3190 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3206 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3222 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3238 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3254 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3270 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3286 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3302 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3318 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3334 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3350 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3366 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3382 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3398 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3414 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3430 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3446 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3462 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3478 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3494 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3510 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3526 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3542 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3558 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3574 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3590 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3606 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3622 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_3638 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_3646 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3670 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3686 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3702 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3718 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3734 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3750 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3766 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3782 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3798 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3814 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3830 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3846 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3862 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3878 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3894 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3910 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3926 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3942 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3958 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3974 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_3990 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4006 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4022 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4038 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4054 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4070 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4086 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4102 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4118 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4134 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4150 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4166 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4182 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_4198 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_4206 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4230 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4246 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4262 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4278 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4294 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4310 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4326 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4342 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4358 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4374 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4390 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4406 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4422 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4438 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4454 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4470 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4486 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4502 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4518 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4534 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4550 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4566 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4582 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4598 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4614 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4630 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4646 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4662 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4678 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4694 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4710 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4726 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4742 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_4758 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_4766 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4790 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4806 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4822 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4838 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4854 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4870 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4886 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4902 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4918 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4934 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4950 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4966 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4982 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_4998 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5014 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5030 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5046 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5062 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5078 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5094 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5110 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5126 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5142 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5158 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5174 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5190 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5206 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5222 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5238 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5254 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5270 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5286 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5302 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_5318 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_5326 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5350 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5366 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5382 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5398 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5414 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5430 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5446 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5462 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5478 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5494 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5510 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5526 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5542 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5558 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5574 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5590 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5606 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5622 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5638 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5654 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5670 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5686 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5702 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5718 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5734 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5750 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5766 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5782 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5798 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5814 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5830 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5846 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5862 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_5878 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_5886 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5910 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5926 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5942 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5958 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5974 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_5990 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6006 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6022 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6038 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6054 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6070 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6086 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6102 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6118 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6134 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6150 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6166 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6182 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6198 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6214 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6230 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6246 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6262 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6278 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6294 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6310 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6326 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6342 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6358 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6374 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6390 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6406 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6422 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_6438 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_6446 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6470 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6486 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6502 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6518 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6534 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6550 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6566 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6582 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6598 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6614 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6630 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6646 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6662 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6678 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6694 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6710 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6726 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6742 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6758 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6774 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6790 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6806 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6822 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6838 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6854 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6870 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6886 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6902 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6918 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6934 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6950 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6966 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_6982 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_6998 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_7006 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7030 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7046 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7062 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7078 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7094 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7110 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7126 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7142 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7158 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7174 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7190 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7206 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7222 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7238 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7254 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7270 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7286 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7302 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7318 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7334 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7350 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7366 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7382 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7398 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7414 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7430 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7446 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7462 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7478 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7494 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7510 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7526 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7542 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_7558 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_7566 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7590 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7606 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7622 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7638 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7654 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7670 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7686 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7702 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7718 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7734 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7750 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7766 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7782 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7798 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7814 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7830 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7846 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7862 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7878 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7894 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7910 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7926 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7942 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7958 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7974 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_7990 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8006 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8022 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8038 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8054 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8070 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8086 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8102 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_8118 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_8126 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8150 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8166 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8182 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8198 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8214 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8230 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8246 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8262 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8278 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8294 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8310 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8326 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8342 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8358 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8374 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8390 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8406 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8422 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8438 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8454 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8470 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8486 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8502 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8518 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8534 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8550 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8566 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8582 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8598 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8614 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8630 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8646 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8662 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_8678 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_8686 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8710 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8726 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8742 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8758 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8774 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8790 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8806 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8822 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8838 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8854 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8870 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8886 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8902 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8918 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8934 ();
 gf180mcu_osu_sc_gp9t3v3__fill_16 FILLER_88_8950 ();
 gf180mcu_osu_sc_gp9t3v3__fill_8 FILLER_88_8966 ();
 gf180mcu_osu_sc_gp9t3v3__fill_2 FILLER_88_8974 ();
 assign o[0] = net1;
 assign o[10] = net11;
 assign o[11] = net12;
 assign o[12] = net13;
 assign o[13] = net14;
 assign o[14] = net15;
 assign o[15] = net16;
 assign o[1] = net2;
 assign o[2] = net3;
 assign o[3] = net4;
 assign o[4] = net5;
 assign o[5] = net6;
 assign o[6] = net7;
 assign o[7] = net8;
 assign o[8] = net9;
 assign o[9] = net10;
endmodule

