magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 453 2102 1094
<< pwell >>
rect -86 -86 2102 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
rect 1468 69 1588 333
rect 1692 69 1812 333
<< mvpmos >>
rect 124 573 224 939
rect 348 573 448 939
rect 572 573 672 939
rect 796 573 896 939
rect 1020 573 1120 939
rect 1244 573 1344 939
rect 1468 573 1568 939
rect 1692 573 1792 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 244 287 348 333
rect 244 147 273 287
rect 319 147 348 287
rect 244 69 348 147
rect 468 287 572 333
rect 468 147 497 287
rect 543 147 572 287
rect 468 69 572 147
rect 692 287 796 333
rect 692 147 721 287
rect 767 147 796 287
rect 692 69 796 147
rect 916 222 1020 333
rect 916 82 945 222
rect 991 82 1020 222
rect 916 69 1020 82
rect 1140 287 1244 333
rect 1140 147 1169 287
rect 1215 147 1244 287
rect 1140 69 1244 147
rect 1364 287 1468 333
rect 1364 147 1393 287
rect 1439 147 1468 287
rect 1364 69 1468 147
rect 1588 287 1692 333
rect 1588 147 1617 287
rect 1663 147 1692 287
rect 1588 69 1692 147
rect 1812 287 1900 333
rect 1812 147 1841 287
rect 1887 147 1900 287
rect 1812 69 1900 147
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 224 861 348 939
rect 224 721 273 861
rect 319 721 348 861
rect 224 573 348 721
rect 448 861 572 939
rect 448 721 477 861
rect 523 721 572 861
rect 448 573 572 721
rect 672 861 796 939
rect 672 721 701 861
rect 747 721 796 861
rect 672 573 796 721
rect 896 861 1020 939
rect 896 721 925 861
rect 971 721 1020 861
rect 896 573 1020 721
rect 1120 861 1244 939
rect 1120 721 1149 861
rect 1195 721 1244 861
rect 1120 573 1244 721
rect 1344 861 1468 939
rect 1344 721 1373 861
rect 1419 721 1468 861
rect 1344 573 1468 721
rect 1568 861 1692 939
rect 1568 721 1597 861
rect 1643 721 1692 861
rect 1568 573 1692 721
rect 1792 861 1880 939
rect 1792 721 1821 861
rect 1867 721 1880 861
rect 1792 573 1880 721
<< mvndiffc >>
rect 49 147 95 287
rect 273 147 319 287
rect 497 147 543 287
rect 721 147 767 287
rect 945 82 991 222
rect 1169 147 1215 287
rect 1393 147 1439 287
rect 1617 147 1663 287
rect 1841 147 1887 287
<< mvpdiffc >>
rect 49 721 95 861
rect 273 721 319 861
rect 477 721 523 861
rect 701 721 747 861
rect 925 721 971 861
rect 1149 721 1195 861
rect 1373 721 1419 861
rect 1597 721 1643 861
rect 1821 721 1867 861
<< polysilicon >>
rect 124 939 224 983
rect 348 939 448 983
rect 572 939 672 983
rect 796 939 896 983
rect 1020 939 1120 983
rect 1244 939 1344 983
rect 1468 939 1568 983
rect 1692 939 1792 983
rect 124 513 224 573
rect 348 513 448 573
rect 572 513 672 573
rect 796 513 896 573
rect 124 512 896 513
rect 1020 513 1120 573
rect 1244 513 1344 573
rect 1468 513 1568 573
rect 1692 513 1792 573
rect 1020 512 1792 513
rect 124 500 1792 512
rect 124 454 137 500
rect 841 454 1072 500
rect 1776 454 1792 500
rect 124 441 1792 454
rect 124 333 244 441
rect 348 333 468 441
rect 572 333 692 441
rect 796 333 916 441
rect 1020 333 1140 441
rect 1244 333 1364 441
rect 1468 333 1588 441
rect 1692 377 1792 441
rect 1692 333 1812 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1468 25 1588 69
rect 1692 25 1812 69
<< polycontact >>
rect 137 454 841 500
rect 1072 454 1776 500
<< metal1 >>
rect 0 918 2016 1098
rect 49 861 95 918
rect 49 710 95 721
rect 273 861 319 872
rect 273 664 319 721
rect 477 861 523 918
rect 477 710 523 721
rect 701 861 747 872
rect 701 664 747 721
rect 925 861 971 918
rect 925 710 971 721
rect 1149 861 1195 872
rect 1149 664 1195 721
rect 1373 861 1419 918
rect 1373 710 1419 721
rect 1597 861 1643 872
rect 1597 664 1643 721
rect 1821 861 1867 918
rect 1821 710 1867 721
rect 273 618 1643 664
rect 126 500 852 529
rect 126 454 137 500
rect 841 454 852 500
rect 126 453 852 454
rect 926 397 1026 618
rect 1072 500 1776 530
rect 1072 443 1776 454
rect 273 351 1663 397
rect 49 287 95 298
rect 49 90 95 147
rect 273 287 319 351
rect 273 136 319 147
rect 497 287 543 298
rect 497 90 543 147
rect 715 287 767 351
rect 715 147 721 287
rect 1169 287 1215 351
rect 715 136 767 147
rect 945 222 991 233
rect 0 82 945 90
rect 1169 136 1215 147
rect 1393 287 1439 298
rect 1393 90 1439 147
rect 1617 287 1663 351
rect 1617 136 1663 147
rect 1841 287 1887 298
rect 1841 90 1887 147
rect 991 82 2016 90
rect 0 -90 2016 82
<< labels >>
flabel metal1 s 126 453 852 529 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 2016 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 1841 233 1887 298 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 1597 664 1643 872 0 FreeSans 200 0 0 0 ZN
port 2 nsew default output
rlabel metal1 s 1072 443 1776 530 1 I
port 1 nsew default input
rlabel metal1 s 1149 664 1195 872 1 ZN
port 2 nsew default output
rlabel metal1 s 701 664 747 872 1 ZN
port 2 nsew default output
rlabel metal1 s 273 664 319 872 1 ZN
port 2 nsew default output
rlabel metal1 s 273 618 1643 664 1 ZN
port 2 nsew default output
rlabel metal1 s 926 397 1026 618 1 ZN
port 2 nsew default output
rlabel metal1 s 273 351 1663 397 1 ZN
port 2 nsew default output
rlabel metal1 s 1617 136 1663 351 1 ZN
port 2 nsew default output
rlabel metal1 s 1169 136 1215 351 1 ZN
port 2 nsew default output
rlabel metal1 s 715 136 767 351 1 ZN
port 2 nsew default output
rlabel metal1 s 273 136 319 351 1 ZN
port 2 nsew default output
rlabel metal1 s 1821 710 1867 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 710 1419 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 710 971 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 710 523 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1393 233 1439 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 233 543 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 233 95 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 90 1887 233 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 233 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 233 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 233 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 233 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2016 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2016 1008
string GDS_END 870024
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 864114
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
