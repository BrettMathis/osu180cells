magic
tech gf180mcuB
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 4480 844
rect 49 629 95 724
rect 467 621 513 724
rect 885 621 931 724
rect 1660 689 1728 724
rect 2409 657 2477 724
rect 2902 657 2970 724
rect 220 403 2094 449
rect 2634 430 2702 577
rect 3170 430 3248 577
rect 220 337 266 403
rect 781 360 1169 403
rect 328 314 694 355
rect 1271 314 1524 357
rect 2634 354 3248 430
rect 328 311 1524 314
rect 328 261 1317 311
rect 328 240 793 261
rect 49 60 95 138
rect 874 60 942 215
rect 2418 60 2488 224
rect 2634 207 2712 354
rect 3180 207 3248 354
rect 3425 546 3471 724
rect 3644 496 3712 678
rect 3879 546 3925 724
rect 4050 496 4169 678
rect 4321 546 4367 724
rect 3644 449 4169 496
rect 4050 274 4169 449
rect 3644 227 4169 274
rect 2912 60 2980 127
rect 3445 60 3491 187
rect 3644 108 3721 227
rect 3888 60 3956 147
rect 4050 130 4169 227
rect 4347 60 4393 187
rect 0 -60 4480 60
<< obsm1 >>
rect 251 563 320 678
rect 670 563 738 678
rect 1144 611 2323 643
rect 2532 623 2811 669
rect 2532 611 2578 623
rect 1144 597 2578 611
rect 2277 565 2578 597
rect 2765 596 2811 623
rect 3063 623 3340 669
rect 3063 596 3109 623
rect 128 551 738 563
rect 128 505 2186 551
rect 128 264 174 505
rect 2140 409 2186 505
rect 2765 550 3109 596
rect 2140 363 2576 409
rect 128 218 251 264
rect 1928 276 2584 317
rect 1577 270 2584 276
rect 1577 265 1996 270
rect 1368 229 1996 265
rect 1368 218 1623 229
rect 1928 218 1996 229
rect 205 154 251 218
rect 205 108 534 154
rect 1144 172 1212 215
rect 1660 172 1728 183
rect 2152 172 2220 215
rect 1144 126 2220 172
rect 2538 152 2584 270
rect 2806 201 3113 247
rect 3294 394 3340 623
rect 3294 348 3972 394
rect 2806 152 2852 201
rect 2538 106 2852 152
rect 3067 152 3113 201
rect 3294 152 3340 348
rect 3067 106 3340 152
<< labels >>
rlabel metal1 s 220 403 2094 449 6 A
port 1 nsew default input
rlabel metal1 s 781 360 1169 403 6 A
port 1 nsew default input
rlabel metal1 s 220 360 266 403 6 A
port 1 nsew default input
rlabel metal1 s 220 337 266 360 6 A
port 1 nsew default input
rlabel metal1 s 1271 355 1524 357 6 B
port 2 nsew default input
rlabel metal1 s 1271 314 1524 355 6 B
port 2 nsew default input
rlabel metal1 s 328 314 694 355 6 B
port 2 nsew default input
rlabel metal1 s 328 311 1524 314 6 B
port 2 nsew default input
rlabel metal1 s 328 261 1317 311 6 B
port 2 nsew default input
rlabel metal1 s 328 240 793 261 6 B
port 2 nsew default input
rlabel metal1 s 3170 430 3248 577 6 CO
port 3 nsew default output
rlabel metal1 s 2634 430 2702 577 6 CO
port 3 nsew default output
rlabel metal1 s 2634 354 3248 430 6 CO
port 3 nsew default output
rlabel metal1 s 3180 207 3248 354 6 CO
port 3 nsew default output
rlabel metal1 s 2634 207 2712 354 6 CO
port 3 nsew default output
rlabel metal1 s 4050 496 4169 678 6 S
port 4 nsew default output
rlabel metal1 s 3644 496 3712 678 6 S
port 4 nsew default output
rlabel metal1 s 3644 449 4169 496 6 S
port 4 nsew default output
rlabel metal1 s 4050 274 4169 449 6 S
port 4 nsew default output
rlabel metal1 s 3644 227 4169 274 6 S
port 4 nsew default output
rlabel metal1 s 4050 130 4169 227 6 S
port 4 nsew default output
rlabel metal1 s 3644 130 3721 227 6 S
port 4 nsew default output
rlabel metal1 s 3644 108 3721 130 6 S
port 4 nsew default output
rlabel metal1 s 0 724 4480 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4321 689 4367 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3879 689 3925 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3425 689 3471 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2902 689 2970 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2409 689 2477 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1660 689 1728 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 885 689 931 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 467 689 513 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 689 95 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4321 657 4367 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3879 657 3925 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3425 657 3471 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2902 657 2970 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2409 657 2477 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 885 657 931 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 467 657 513 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 657 95 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4321 629 4367 657 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3879 629 3925 657 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3425 629 3471 657 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 885 629 931 657 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 467 629 513 657 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 629 95 657 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4321 621 4367 629 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3879 621 3925 629 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3425 621 3471 629 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 885 621 931 629 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 467 621 513 629 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4321 546 4367 621 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3879 546 3925 621 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3425 546 3471 621 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2418 215 2488 224 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2418 187 2488 215 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 874 187 942 215 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4347 147 4393 187 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3445 147 3491 187 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2418 147 2488 187 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 874 147 942 187 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4347 138 4393 147 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3888 138 3956 147 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3445 138 3491 147 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2418 138 2488 147 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 874 138 942 147 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4347 127 4393 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3888 127 3956 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3445 127 3491 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2418 127 2488 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 874 127 942 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 127 95 138 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 4347 60 4393 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3888 60 3956 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3445 60 3491 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2912 60 2980 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2418 60 2488 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 874 60 942 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4480 60 8 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4480 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1185356
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1176828
<< end >>
