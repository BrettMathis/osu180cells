magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< metal1 >>
rect 0 724 448 844
rect 353 498 399 724
rect 49 60 95 219
rect 0 -60 448 60
<< obsm1 >>
rect 49 311 95 678
rect 146 392 399 438
rect 49 265 304 311
rect 353 106 399 392
<< labels >>
rlabel metal1 s 0 724 448 844 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 498 399 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 49 60 95 219 6 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 448 60 8 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 784
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1134414
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1132262
<< end >>
