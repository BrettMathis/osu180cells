magic
tech gf180mcuC
magscale 1 10
timestamp 1669390400
<< nwell >>
rect -86 352 7030 870
<< pwell >>
rect -86 -86 7030 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 1916 68 2036 232
rect 2140 68 2260 232
rect 2364 68 2484 232
rect 2588 68 2708 232
rect 2812 68 2932 232
rect 3036 68 3156 232
rect 3260 68 3380 232
rect 3484 68 3604 232
rect 3708 68 3828 232
rect 3932 68 4052 232
rect 4156 68 4276 232
rect 4380 68 4500 232
rect 4604 68 4724 232
rect 4828 68 4948 232
rect 5052 68 5172 232
rect 5276 68 5396 232
rect 5500 68 5620 232
rect 5724 68 5844 232
rect 5948 68 6068 232
rect 6172 68 6292 232
rect 6396 68 6516 232
rect 6620 68 6740 232
<< mvpmos >>
rect 124 472 224 716
rect 348 472 448 716
rect 572 472 672 716
rect 796 472 896 716
rect 1020 472 1120 716
rect 1244 472 1344 716
rect 1468 472 1568 716
rect 1692 472 1792 716
rect 1916 472 2016 716
rect 2140 472 2240 716
rect 2364 472 2464 716
rect 2588 472 2688 716
rect 2812 472 2912 716
rect 3036 472 3136 716
rect 3260 472 3360 716
rect 3484 472 3584 716
rect 3708 472 3808 716
rect 3932 472 4032 716
rect 4156 472 4256 716
rect 4380 472 4480 716
rect 4604 472 4704 716
rect 4828 472 4928 716
rect 5052 472 5152 716
rect 5276 472 5376 716
rect 5500 472 5600 716
rect 5724 472 5824 716
rect 5948 472 6048 716
rect 6172 472 6272 716
rect 6396 472 6496 716
rect 6620 472 6720 716
<< mvndiff >>
rect 36 192 124 232
rect 36 146 49 192
rect 95 146 124 192
rect 36 68 124 146
rect 244 192 348 232
rect 244 146 273 192
rect 319 146 348 192
rect 244 68 348 146
rect 468 181 572 232
rect 468 135 497 181
rect 543 135 572 181
rect 468 68 572 135
rect 692 192 796 232
rect 692 146 721 192
rect 767 146 796 192
rect 692 68 796 146
rect 916 181 1020 232
rect 916 135 945 181
rect 991 135 1020 181
rect 916 68 1020 135
rect 1140 192 1244 232
rect 1140 146 1169 192
rect 1215 146 1244 192
rect 1140 68 1244 146
rect 1364 181 1468 232
rect 1364 135 1393 181
rect 1439 135 1468 181
rect 1364 68 1468 135
rect 1588 192 1692 232
rect 1588 146 1617 192
rect 1663 146 1692 192
rect 1588 68 1692 146
rect 1812 181 1916 232
rect 1812 135 1841 181
rect 1887 135 1916 181
rect 1812 68 1916 135
rect 2036 192 2140 232
rect 2036 146 2065 192
rect 2111 146 2140 192
rect 2036 68 2140 146
rect 2260 181 2364 232
rect 2260 135 2289 181
rect 2335 135 2364 181
rect 2260 68 2364 135
rect 2484 192 2588 232
rect 2484 146 2513 192
rect 2559 146 2588 192
rect 2484 68 2588 146
rect 2708 127 2812 232
rect 2708 81 2737 127
rect 2783 81 2812 127
rect 2708 68 2812 81
rect 2932 192 3036 232
rect 2932 146 2961 192
rect 3007 146 3036 192
rect 2932 68 3036 146
rect 3156 127 3260 232
rect 3156 81 3185 127
rect 3231 81 3260 127
rect 3156 68 3260 81
rect 3380 192 3484 232
rect 3380 146 3409 192
rect 3455 146 3484 192
rect 3380 68 3484 146
rect 3604 127 3708 232
rect 3604 81 3633 127
rect 3679 81 3708 127
rect 3604 68 3708 81
rect 3828 192 3932 232
rect 3828 146 3857 192
rect 3903 146 3932 192
rect 3828 68 3932 146
rect 4052 127 4156 232
rect 4052 81 4081 127
rect 4127 81 4156 127
rect 4052 68 4156 81
rect 4276 192 4380 232
rect 4276 146 4305 192
rect 4351 146 4380 192
rect 4276 68 4380 146
rect 4500 127 4604 232
rect 4500 81 4529 127
rect 4575 81 4604 127
rect 4500 68 4604 81
rect 4724 192 4828 232
rect 4724 146 4753 192
rect 4799 146 4828 192
rect 4724 68 4828 146
rect 4948 127 5052 232
rect 4948 81 4977 127
rect 5023 81 5052 127
rect 4948 68 5052 81
rect 5172 192 5276 232
rect 5172 146 5201 192
rect 5247 146 5276 192
rect 5172 68 5276 146
rect 5396 127 5500 232
rect 5396 81 5425 127
rect 5471 81 5500 127
rect 5396 68 5500 81
rect 5620 192 5724 232
rect 5620 146 5649 192
rect 5695 146 5724 192
rect 5620 68 5724 146
rect 5844 127 5948 232
rect 5844 81 5873 127
rect 5919 81 5948 127
rect 5844 68 5948 81
rect 6068 192 6172 232
rect 6068 146 6097 192
rect 6143 146 6172 192
rect 6068 68 6172 146
rect 6292 127 6396 232
rect 6292 81 6321 127
rect 6367 81 6396 127
rect 6292 68 6396 81
rect 6516 192 6620 232
rect 6516 146 6545 192
rect 6591 146 6620 192
rect 6516 68 6620 146
rect 6740 192 6828 232
rect 6740 146 6769 192
rect 6815 146 6828 192
rect 6740 68 6828 146
<< mvpdiff >>
rect 36 665 124 716
rect 36 525 49 665
rect 95 525 124 665
rect 36 472 124 525
rect 224 665 348 716
rect 224 525 273 665
rect 319 525 348 665
rect 224 472 348 525
rect 448 665 572 716
rect 448 619 477 665
rect 523 619 572 665
rect 448 472 572 619
rect 672 665 796 716
rect 672 525 701 665
rect 747 525 796 665
rect 672 472 796 525
rect 896 665 1020 716
rect 896 619 925 665
rect 971 619 1020 665
rect 896 472 1020 619
rect 1120 665 1244 716
rect 1120 525 1149 665
rect 1195 525 1244 665
rect 1120 472 1244 525
rect 1344 665 1468 716
rect 1344 619 1373 665
rect 1419 619 1468 665
rect 1344 472 1468 619
rect 1568 665 1692 716
rect 1568 525 1597 665
rect 1643 525 1692 665
rect 1568 472 1692 525
rect 1792 665 1916 716
rect 1792 619 1821 665
rect 1867 619 1916 665
rect 1792 472 1916 619
rect 2016 665 2140 716
rect 2016 525 2045 665
rect 2091 525 2140 665
rect 2016 472 2140 525
rect 2240 665 2364 716
rect 2240 525 2269 665
rect 2315 525 2364 665
rect 2240 472 2364 525
rect 2464 665 2588 716
rect 2464 525 2513 665
rect 2559 525 2588 665
rect 2464 472 2588 525
rect 2688 703 2812 716
rect 2688 657 2717 703
rect 2763 657 2812 703
rect 2688 472 2812 657
rect 2912 665 3036 716
rect 2912 525 2941 665
rect 2987 525 3036 665
rect 2912 472 3036 525
rect 3136 703 3260 716
rect 3136 657 3165 703
rect 3211 657 3260 703
rect 3136 472 3260 657
rect 3360 665 3484 716
rect 3360 525 3389 665
rect 3435 525 3484 665
rect 3360 472 3484 525
rect 3584 703 3708 716
rect 3584 657 3613 703
rect 3659 657 3708 703
rect 3584 472 3708 657
rect 3808 665 3932 716
rect 3808 525 3837 665
rect 3883 525 3932 665
rect 3808 472 3932 525
rect 4032 703 4156 716
rect 4032 657 4061 703
rect 4107 657 4156 703
rect 4032 472 4156 657
rect 4256 665 4380 716
rect 4256 525 4285 665
rect 4331 525 4380 665
rect 4256 472 4380 525
rect 4480 703 4604 716
rect 4480 657 4509 703
rect 4555 657 4604 703
rect 4480 472 4604 657
rect 4704 665 4828 716
rect 4704 525 4733 665
rect 4779 525 4828 665
rect 4704 472 4828 525
rect 4928 703 5052 716
rect 4928 657 4957 703
rect 5003 657 5052 703
rect 4928 472 5052 657
rect 5152 665 5276 716
rect 5152 525 5181 665
rect 5227 525 5276 665
rect 5152 472 5276 525
rect 5376 703 5500 716
rect 5376 657 5405 703
rect 5451 657 5500 703
rect 5376 472 5500 657
rect 5600 665 5724 716
rect 5600 525 5629 665
rect 5675 525 5724 665
rect 5600 472 5724 525
rect 5824 703 5948 716
rect 5824 657 5853 703
rect 5899 657 5948 703
rect 5824 472 5948 657
rect 6048 665 6172 716
rect 6048 525 6077 665
rect 6123 525 6172 665
rect 6048 472 6172 525
rect 6272 703 6396 716
rect 6272 657 6301 703
rect 6347 657 6396 703
rect 6272 472 6396 657
rect 6496 665 6620 716
rect 6496 525 6525 665
rect 6571 525 6620 665
rect 6496 472 6620 525
rect 6720 665 6808 716
rect 6720 525 6749 665
rect 6795 525 6808 665
rect 6720 472 6808 525
<< mvndiffc >>
rect 49 146 95 192
rect 273 146 319 192
rect 497 135 543 181
rect 721 146 767 192
rect 945 135 991 181
rect 1169 146 1215 192
rect 1393 135 1439 181
rect 1617 146 1663 192
rect 1841 135 1887 181
rect 2065 146 2111 192
rect 2289 135 2335 181
rect 2513 146 2559 192
rect 2737 81 2783 127
rect 2961 146 3007 192
rect 3185 81 3231 127
rect 3409 146 3455 192
rect 3633 81 3679 127
rect 3857 146 3903 192
rect 4081 81 4127 127
rect 4305 146 4351 192
rect 4529 81 4575 127
rect 4753 146 4799 192
rect 4977 81 5023 127
rect 5201 146 5247 192
rect 5425 81 5471 127
rect 5649 146 5695 192
rect 5873 81 5919 127
rect 6097 146 6143 192
rect 6321 81 6367 127
rect 6545 146 6591 192
rect 6769 146 6815 192
<< mvpdiffc >>
rect 49 525 95 665
rect 273 525 319 665
rect 477 619 523 665
rect 701 525 747 665
rect 925 619 971 665
rect 1149 525 1195 665
rect 1373 619 1419 665
rect 1597 525 1643 665
rect 1821 619 1867 665
rect 2045 525 2091 665
rect 2269 525 2315 665
rect 2513 525 2559 665
rect 2717 657 2763 703
rect 2941 525 2987 665
rect 3165 657 3211 703
rect 3389 525 3435 665
rect 3613 657 3659 703
rect 3837 525 3883 665
rect 4061 657 4107 703
rect 4285 525 4331 665
rect 4509 657 4555 703
rect 4733 525 4779 665
rect 4957 657 5003 703
rect 5181 525 5227 665
rect 5405 657 5451 703
rect 5629 525 5675 665
rect 5853 657 5899 703
rect 6077 525 6123 665
rect 6301 657 6347 703
rect 6525 525 6571 665
rect 6749 525 6795 665
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 572 716 672 760
rect 796 716 896 760
rect 1020 716 1120 760
rect 1244 716 1344 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1916 716 2016 760
rect 2140 716 2240 760
rect 2364 716 2464 760
rect 2588 716 2688 760
rect 2812 716 2912 760
rect 3036 716 3136 760
rect 3260 716 3360 760
rect 3484 716 3584 760
rect 3708 716 3808 760
rect 3932 716 4032 760
rect 4156 716 4256 760
rect 4380 716 4480 760
rect 4604 716 4704 760
rect 4828 716 4928 760
rect 5052 716 5152 760
rect 5276 716 5376 760
rect 5500 716 5600 760
rect 5724 716 5824 760
rect 5948 716 6048 760
rect 6172 716 6272 760
rect 6396 716 6496 760
rect 6620 716 6720 760
rect 124 407 224 472
rect 348 407 448 472
rect 572 407 672 472
rect 796 407 896 472
rect 1020 407 1120 472
rect 1244 407 1344 472
rect 1468 407 1568 472
rect 1692 407 1792 472
rect 1916 407 2016 472
rect 124 394 2016 407
rect 2140 394 2240 472
rect 124 348 137 394
rect 1969 350 2240 394
rect 1969 348 2036 350
rect 124 335 2036 348
rect 124 232 244 335
rect 348 232 468 335
rect 572 232 692 335
rect 796 232 916 335
rect 1020 232 1140 335
rect 1244 232 1364 335
rect 1468 232 1588 335
rect 1692 232 1812 335
rect 1916 232 2036 335
rect 2140 288 2240 350
rect 2364 407 2464 472
rect 2588 407 2688 472
rect 2812 407 2912 472
rect 3036 407 3136 472
rect 3260 407 3360 472
rect 3484 407 3584 472
rect 3708 407 3808 472
rect 3932 407 4032 472
rect 4156 407 4256 472
rect 4380 407 4480 472
rect 4604 407 4704 472
rect 4828 407 4928 472
rect 5052 407 5152 472
rect 5276 407 5376 472
rect 5500 407 5600 472
rect 5724 407 5824 472
rect 5948 407 6048 472
rect 6172 407 6272 472
rect 6396 407 6496 472
rect 6620 407 6720 472
rect 2364 394 6720 407
rect 2364 348 2377 394
rect 4303 348 4747 394
rect 6673 348 6720 394
rect 2364 335 6720 348
rect 2140 232 2260 288
rect 2364 232 2484 335
rect 2588 232 2708 335
rect 2812 232 2932 335
rect 3036 232 3156 335
rect 3260 232 3380 335
rect 3484 232 3604 335
rect 3708 232 3828 335
rect 3932 232 4052 335
rect 4156 232 4276 335
rect 4380 232 4500 335
rect 4604 232 4724 335
rect 4828 232 4948 335
rect 5052 232 5172 335
rect 5276 232 5396 335
rect 5500 232 5620 335
rect 5724 232 5844 335
rect 5948 232 6068 335
rect 6172 232 6292 335
rect 6396 232 6516 335
rect 6620 288 6720 335
rect 6620 232 6740 288
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 1916 24 2036 68
rect 2140 24 2260 68
rect 2364 24 2484 68
rect 2588 24 2708 68
rect 2812 24 2932 68
rect 3036 24 3156 68
rect 3260 24 3380 68
rect 3484 24 3604 68
rect 3708 24 3828 68
rect 3932 24 4052 68
rect 4156 24 4276 68
rect 4380 24 4500 68
rect 4604 24 4724 68
rect 4828 24 4948 68
rect 5052 24 5172 68
rect 5276 24 5396 68
rect 5500 24 5620 68
rect 5724 24 5844 68
rect 5948 24 6068 68
rect 6172 24 6292 68
rect 6396 24 6516 68
rect 6620 24 6740 68
<< polycontact >>
rect 137 348 1969 394
rect 2377 348 4303 394
rect 4747 348 6673 394
<< metal1 >>
rect 0 724 6944 844
rect 49 665 95 724
rect 49 506 95 525
rect 273 665 319 676
rect 477 665 523 724
rect 477 600 523 619
rect 701 665 747 676
rect 319 525 701 552
rect 925 665 971 724
rect 925 600 971 619
rect 1149 665 1195 676
rect 747 525 1149 552
rect 1373 665 1419 724
rect 1373 600 1419 619
rect 1597 665 1643 676
rect 1195 525 1597 552
rect 1821 665 1867 724
rect 1821 600 1867 619
rect 2045 665 2136 676
rect 1643 525 2045 552
rect 2091 525 2136 665
rect 273 506 2136 525
rect 2269 665 2315 724
rect 2717 703 2763 724
rect 2269 506 2315 525
rect 2513 665 2559 676
rect 3165 703 3211 724
rect 2717 646 2763 657
rect 2941 665 2987 676
rect 2559 525 2941 600
rect 3613 703 3659 724
rect 3165 646 3211 657
rect 3389 665 3435 676
rect 2987 525 3389 600
rect 4061 703 4107 724
rect 3613 646 3659 657
rect 3837 665 3883 676
rect 3435 525 3837 600
rect 4509 703 4555 724
rect 4061 646 4107 657
rect 4285 665 4331 676
rect 3883 525 4285 600
rect 4957 703 5003 724
rect 4509 646 4555 657
rect 4733 665 4779 676
rect 4331 525 4733 600
rect 5405 703 5451 724
rect 4957 646 5003 657
rect 5181 665 5227 676
rect 4779 525 5181 600
rect 5853 703 5899 724
rect 5405 646 5451 657
rect 5629 665 5675 676
rect 5227 525 5629 600
rect 6301 703 6347 724
rect 5853 646 5899 657
rect 6077 665 6123 676
rect 5675 525 6077 600
rect 6301 646 6347 657
rect 6525 665 6571 676
rect 6123 525 6525 600
rect 126 394 1980 430
rect 126 348 137 394
rect 1969 348 1980 394
rect 2045 394 2136 506
rect 2513 454 6571 525
rect 6749 665 6795 724
rect 6749 506 6795 525
rect 2045 348 2377 394
rect 4303 348 4314 394
rect 2045 284 2136 348
rect 4446 302 4626 454
rect 4736 348 4747 394
rect 6673 348 6720 394
rect 273 238 2136 284
rect 49 192 95 232
rect 49 60 95 146
rect 273 192 319 238
rect 721 192 767 238
rect 1169 192 1215 238
rect 1617 192 1663 238
rect 2065 192 2136 238
rect 2513 192 6591 302
rect 273 135 319 146
rect 497 181 543 192
rect 721 135 767 146
rect 945 181 991 192
rect 1169 135 1215 146
rect 1393 181 1439 192
rect 1617 135 1663 146
rect 1841 181 1887 192
rect 2111 146 2136 192
rect 2065 135 2136 146
rect 2289 181 2335 192
rect 2559 173 2961 192
rect 2559 146 2565 173
rect 2513 135 2565 146
rect 3007 173 3409 192
rect 2961 135 3007 146
rect 3455 173 3857 192
rect 3409 135 3455 146
rect 3903 173 4305 192
rect 3857 135 3903 146
rect 4351 173 4753 192
rect 4305 135 4351 146
rect 4799 173 5201 192
rect 4753 135 4799 146
rect 5247 173 5649 192
rect 5201 135 5247 146
rect 5695 173 6097 192
rect 5649 135 5695 146
rect 6143 173 6545 192
rect 6097 135 6143 146
rect 6545 135 6591 146
rect 6769 192 6815 232
rect 497 60 543 135
rect 945 60 991 135
rect 1393 60 1439 135
rect 1841 60 1887 135
rect 2289 60 2335 135
rect 2726 81 2737 127
rect 2783 81 2794 127
rect 2726 60 2794 81
rect 3174 81 3185 127
rect 3231 81 3242 127
rect 3174 60 3242 81
rect 3622 81 3633 127
rect 3679 81 3690 127
rect 3622 60 3690 81
rect 4070 81 4081 127
rect 4127 81 4138 127
rect 4070 60 4138 81
rect 4518 81 4529 127
rect 4575 81 4586 127
rect 4518 60 4586 81
rect 4966 81 4977 127
rect 5023 81 5034 127
rect 4966 60 5034 81
rect 5414 81 5425 127
rect 5471 81 5482 127
rect 5414 60 5482 81
rect 5862 81 5873 127
rect 5919 81 5930 127
rect 5862 60 5930 81
rect 6310 81 6321 127
rect 6367 81 6378 127
rect 6310 60 6378 81
rect 6769 60 6815 146
rect 0 -60 6944 60
<< labels >>
flabel metal1 s 0 724 6944 844 0 FreeSans 600 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 6769 192 6815 232 0 FreeSans 600 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 6525 600 6571 676 0 FreeSans 600 0 0 0 Z
port 2 nsew default output
flabel metal1 s 126 348 1980 430 0 FreeSans 600 0 0 0 I
port 1 nsew default input
rlabel metal1 s 6077 600 6123 676 1 Z
port 2 nsew default output
rlabel metal1 s 5629 600 5675 676 1 Z
port 2 nsew default output
rlabel metal1 s 5181 600 5227 676 1 Z
port 2 nsew default output
rlabel metal1 s 4733 600 4779 676 1 Z
port 2 nsew default output
rlabel metal1 s 4285 600 4331 676 1 Z
port 2 nsew default output
rlabel metal1 s 3837 600 3883 676 1 Z
port 2 nsew default output
rlabel metal1 s 3389 600 3435 676 1 Z
port 2 nsew default output
rlabel metal1 s 2941 600 2987 676 1 Z
port 2 nsew default output
rlabel metal1 s 2513 600 2559 676 1 Z
port 2 nsew default output
rlabel metal1 s 2513 454 6571 600 1 Z
port 2 nsew default output
rlabel metal1 s 4446 302 4626 454 1 Z
port 2 nsew default output
rlabel metal1 s 2513 173 6591 302 1 Z
port 2 nsew default output
rlabel metal1 s 6545 135 6591 173 1 Z
port 2 nsew default output
rlabel metal1 s 6097 135 6143 173 1 Z
port 2 nsew default output
rlabel metal1 s 5649 135 5695 173 1 Z
port 2 nsew default output
rlabel metal1 s 5201 135 5247 173 1 Z
port 2 nsew default output
rlabel metal1 s 4753 135 4799 173 1 Z
port 2 nsew default output
rlabel metal1 s 4305 135 4351 173 1 Z
port 2 nsew default output
rlabel metal1 s 3857 135 3903 173 1 Z
port 2 nsew default output
rlabel metal1 s 3409 135 3455 173 1 Z
port 2 nsew default output
rlabel metal1 s 2961 135 3007 173 1 Z
port 2 nsew default output
rlabel metal1 s 2513 135 2565 173 1 Z
port 2 nsew default output
rlabel metal1 s 6749 646 6795 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6301 646 6347 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5853 646 5899 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 646 5451 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4957 646 5003 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 646 4555 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4061 646 4107 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 646 3659 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 646 3211 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 646 2763 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 646 2315 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 646 1867 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 646 1419 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 646 971 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 646 523 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 646 95 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6749 600 6795 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 600 2315 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 600 1867 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 600 1419 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 600 971 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 600 523 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 600 95 646 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6749 506 6795 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 506 2315 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 600 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 192 95 232 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6769 127 6815 192 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 127 2335 192 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 127 1887 192 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 127 1439 192 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 127 991 192 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 127 543 192 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 127 95 192 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6769 60 6815 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6310 60 6378 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5862 60 5930 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5414 60 5482 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4966 60 5034 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4518 60 4586 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 60 2335 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 60 1887 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 60 1439 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 6944 60 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6944 784
string GDS_END 1359712
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1345148
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
